��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�6�!�~�\@NQzB5�1�kR8�W��7�����e6� �����ْ����5�}܇��M� f�/�_�p���Y۪�^�ow��PS�*'��,e�/�W^j��������ք��ݜQRiZ�-
�}u�d�|"4�����fTD~e{�I��ks�W�oKG��]��6Du������V���r@�Wcle5�t��"��a�ǎ����"b:ٯ��O�A���k���֩y
�^P��}cC5	,R�W)��ɑ"�C��Wh9U�sɕ�B{�T��'���Ч�k/Ƭ��7�kֳ�q��	�c8Y�&s�mCM���lZ�~>�f7@��(�a�JL/��������Ly���C�2g�& ;���ս�\w���Hu���4J4Y���!P*Z_|޼��1xA�/���m�������/&���Cʿ(
��,@�d܈�K����~?8�d���s�s��c�8܂��l���SX��G2�`�<Tt5iP&JP�2�8|�1*�)юa��А�t������p���������7?}�s�{��־���l����M}�)� _
�o��&pPW>���X+R�T��<�V������4�\-N�����U�g H3$#6
�q�֕�,Wz}��E��ۅ��Zdc��(���f�6 "4����a�O̀�R�mrM��?��Cgh��7L�����43K�ե��Ƈ���3ylc���}�Ū�`O��b��R�|t�����.���!�F#�0�}.*:"���|�����Z:E�\�d�I�\Q0����v�֯w�j����Ć,{�+b�Q~�X0�h�(D���p;蜁�!p+~MP�O��X#-t��f}Ɏo��`R>V>�����^��]W�X$�7ˀ����KҚڥ�}��7�����*�דyRQ��#[�H"Q+���A�ÿD{�@�
��LH=֜B_�,g�B@P�S*�[f�y�1�+b������N��l�e(<B��R����(�yu�)��?����O]��EW���(jʄ��t��G���K��EӮf��_�E��vQO�e�ƻ��mՀe��L$�$�=���dr�:�Ru��lJ�]��Ʃ+Q5�S|�A0L����c��/���)NOo[.��6���/U�n��M6-^F��RQ8Xu�:�ɧ����XG%�Փ�xV���xo`5,�`ϻ���#�G���ە˧�yQrG�?���&��A%1�"cu_	�Yէg7?�����E@<{���F��3y��������Jr�]�:UyrP��m����y�C�n�%�M�������}��|�a֪��ݾ�7�K�Δ1���2S
XύsO<�1�?��M͢�
B{�����οLқq	�s��F��C��N\H�gj��'%[�:U.&��x�I7�9�&��%M�|~-!墸��h����c�Z	m������ Kr�oS��n�bP��F3Ӛy
��������ێ����pe@#����|\�+K@�HU��G�9�K� ��r�󧴺���@���E���T�7����<�/xz�����a<<6p�:���+��]i�"�F�����c?^ Xb3�/�
�S`�v���Eץ	<�	٨�[V4t�E���w$���ƙv1��m+d�<��	����b.����^wY�$�y<���g�F����W�]��~-r�L�ϴ>���-X>�@C�J36�j�RYT�8���H'����!(Е�e�f5����Z2��#엁���2�Xa���ϹL3�ݿ:a�bc��%�HbF<UP$����[	��|#/v���ě�����S1�7�i��Uz2D�jpQ���	۲G^�ddo�&����٨�h-�IvE�'�5�>J�՞���q-�h1��3�M�3m8u�G�(��ƽ��Éί�x�c�t�Qu�2i���<������O>�p!a�x~�٨p$"���&4,�w�e�[X�'� ����s�p[A���nW��Ib�\s-2�;zX3�p�	�Ou��s�\al��Aکφoy�GY\��ֲs@7��M	��Y�W,G������˅�{<�xw�����t�\H�I��.mcn�Ť��T��[ї�m���%{1ez������k[31;[ yƣy'�Z�% C�QK1�2���t��?��C��ԇ��߻�p�������r�������:���Ӡ�-�p��\�/��A{����A{qŽ����%����n=�NH@�5큲H�oٗ��@gb+̱?gI{��̅Q��3��'����lT�h�	ʿ�-����{Gp��u�k�y��J�p���F>�8�\h|� !׮$X��7>���積Dk��Y�&8�O��HO2����{�9�:@*��wdg!��K`����'ws!�٠|�T��T����f�l�or���%��";Q��	I��\<���9����m4�����"���4ˀ����A̓�b�T@�&s# ����4�E�nZ���>����.�0B*C�q9���a��Eʄ%T{�cR��il\Ԛ���dt���)�� 3k��'0���Ndݶ��}��f������Z�q*��$��j-�&F��iD��*�(�ٻ�X�aʅJ%��P���� �n!����5����'E�Eы�ՋMИ��Ɇ�A�HQ�76�/�%�#v���2=�'�)F¤�pQ�����4~s�b�Ҩ�Aw���*�=z�Տ2��롉ڴ�e�7�Bc�]��uK7_�����r#i�j�tL
���l8�����ܹU�N����S�]Df�	��r���!]�W�ӂ���') �kN4�>��j[~.�`�a��p�r�u{�\�O�>�t��qP����,Z�7ՄXyU��yRyC�F�y��1$�7�vY=��KK��4g6.�;�'��f�=�'��@�~Me�X���{v<r�%��̓v���	sI����.+���o��dޠ� �[�c$��;��j����>N\c��(ּԸ� �����PDO�G���(���CL��.E|�_50"0 �\N����]�a0vc���1���)\�k��������BtD������	)��T��&��/�V6+%"Չ~�*��r�����s���y� K��~�р��vM��N����{��X��M΄�q}h��al^I-��Ou�?�����^�&>��]EՅ"�������TI�+V?fVY�b
��M��V�sd���C��<����CmF�����/#�\�I$�@y�<�*ϛ*���6I�hj�-�(�@�%���m��a�wj�N�3%Z�$��N�̬tz�2�2�NZ�3hݷm���p��eaI�������?����im�Q��G���K[L܁r���W˸LɗP�a����f���8�0m��ڹ]�Q���f�a'�k�_�
l�6�fQa�Ƨ�����s��ʝ�GKuw�H'e��GQ<G�H��t�ڈ�j�h�Ӿ4����xjYD����y����JS5{�
�g���.��)�PQ��3Ǥɑ������m`��_cBI"����b�'�B_��g+���v����'��M��
�[r��}D1G�����~>�[&��nTq�:�RV�bM۾�j�]q̲�ԍ���JĢ����1!j�j�����������:��Al��OOc�]�$�/�ί��6*��+�[���ƒF�t��D)���Sstܢ(�����>����z~Ğ�R_�뽾Z�h܆`7�Q����O�T*5����;g֍p	[-�c$Bβ$v.\KЄ�p!�p�;!9]��_�dt+�Ǩ�����&��6��U�z�L?�)I�+/΃�"�m���k���~�zl��Ćx��ۥ���K1��cT�=֤*�b�qYD����t Ki�B�z�đ�wh�tz�*<�Ѿ�'+���i�a�+�yKv�C��:�ȟ�q}ۇu9Ym�R��$-r�|a���jqF�q@��2<] �vr�'��r׻�v��H��~����8On�b ��:-��3���=z��r3Y�htQD��!Ɏ���x�y=EJSkq�7��шS�!�����^��sڿ)�V+��?����l��W~:3+N\N�mCn\G|	FJ�N-��	�����cN;k�-l���]%ė������gh�J3������ԫ~����$�*��u�zp�Ip�[���i[�/�=,f�~쓐����7˷x� g�c��n�t���H3.�]�R�Y�k/�G�%%�W���! �]��Ƣ���ȴH%JI��^��f϶d�n�.���D�5!I�Z���H������^?�<�'�&�I�&���jo�&Tl���C�V�GA�Rz��h�*먞ӽ��;�Told�U��N�vR�V�5�N���/ysY}�)i&nMS�9(�}�IRM�
��.�r���Bݭ��p^#ĥ�t���,�ڈI���;�
g�{�9Zif��r�)+t�Af\�M
O�y�D|D[6�Sܕ�����aw8�(�G\��"���o�°�Rr�Pvxl�ɝ��\s�e˦�K`���W��6�t���\�;�zg�Bj;���	�
�iO�	�%����Ci�%\�����߲0�&Mw���e�Rr{�߰�U�dL�zs ��d,�CZ���qW|�.Zߔ� vgd�)�Z�rm�s�i���~�a��!�N�GW�e�j��Nr���矻En����v��g�⺒á�
-7�F����ē��̀���.��I�2j
Z�84��L)�OCp�:�E�X���j�A0{��G�C���Od�G!w��'���N�����:	�]]h)��o"�o���"YU�N؟L�w1P����;��89*1�����q��x�^~�ٱ['tL]/�Z�c�H���Өn���7�h�n���Cp05���{t�#�9��)V*���5$�����fQU7{�-��3P�+��잴����'�9]�I{��S�$��dޑT�� ��]}��GR�#��ؖ�~�Q^�D�೙<+��XF��ԗ�1��Ĥ���vg�U/�Ɖ�/},��U7���)1,�Q�C�������8,�gb��56ԝC%�&��o*`�e���\B>n�J	��G�$i�}C��M�=C��!r�'�V�ڎ\�t�)��������=�4e;�� 0(�W�k��\kb9n>��]x$������N�O ]�1c$�>���7w���8�#��w��Ѿ�e1�|��އ���I�B���u�Z{��^�mS���g�A@�����/hI|^�$)�@\� �Z���$��i���Lج�;R�5��̽���Y�1���p)ڄF���#�H�P�d��t���N�T�Nb!�����U����_�F�`c�di��$�Հ�k�^�Qq�����)M�ũ�y|}�yfs�)������Brz�#�W���\z�5���Y)]^�'�:д�(C�� 1��	TU��+���b(��-o�[���O�r�^D�\}�?k�
�>�a�g)b����x�<�F;�5'�~,vd7�7/Z0�Y�>u �ݢj�z�P���0�Vmc���j��Wk�A̡m��=�F�oـ;�$��� 4�It�o4��Ib���!���B�:8,�{5������`����\��
8p@^mP�9S
�yX�;-�$�Xk���QN�	^�Z����=Ԓ:����f��Ί\�%�����BΠ��i��[_>�����vu��c�j�YB�LƧ���2i�S?���'���uG��f�؜�d�<�<���\X����.�:s�5_N�����#������%�4�o�����&p�@ȥ�[��P�D�S���f
=�5ط�ؼ�W��2�E�t�4GflK
Q��B��^-��_���h{���dc~$�ފ��#��tҠj[iy
�#�{?�Ni(�iM1���2��9���b����2o���ˈnAI�	|��Ƕ�4N�_?]��פ�<�eL������Ӻ��`�xޟ����M5&�Pbnn�5��UA�)Qdؼz��h��U��>���P��s����24/�cF+[��j��@��ā��B�q̺_�A*L Fr-6�Ѝ��3��4¥B�`u�&�{���2�W����M�8/a`�������f�v���
}-�����Z㨜zӷ�"Xs��_z�)2CG�� ���U &�l�c��Ob��׈ڃ�pK���:;#y����;��Æ��(��'^�2;Em�#��$�H̫� ['J� U�x��ٱ�n1�a�d0Iv[7NT���qno5Px�y�9�ӂ�\�������*<�q|O���`�%�gh���������y(������qi�j����r�Dua�T3Ղ
_<=�5g����
���M˦&�\�����2�l
tJ�GqC7�e�w�}is�7߭�Ro��#
�1����>�3Q�곭l쨁�-�3ϴΣv�WؤF<��C{�����p���k��؅~*p�;��k�(DK�'d�_��֎��eS����	g=|R���S��ɟh���v�X�X�g��|���&8e��]�k������>���~��0�R. ��9ѿ�w�̺^�7���,�5�z�?���:KAn��
�����W�:P
a�j�V��#h�Y�E��{�[հ"~��Ѵ�7l����V�Ԁ,�?c�7�<+�Åh�$��4�Ru=�,5.���E�7Z*���i"d���u�W �!�mg��U���d~����1<��\4M��&����夃�4�|�i��=��C�U?�)ڱX~I���v��sCOC�����B� '���ke���#C8��n��g�^'w_v��] ���¢[F���D�I7b����S����9�Ĩ������w���fv*��yw;�Z[�7,%0->}T��&�5iSD�JF�3H"����I~�s3��[z6�9N�\"n��z�xq&(X�7�K]p�?,c^}+�F�4/fѼ����D�7��O���:��ܗ�ui�������+�W�5+�Y�~�A��TZ��.k%�V��U�h6�V�|z��j\��NU�aS]�Q�J�7ڙR���t+&V�i��]LP�0oȘ�������3}�>ݸq�����U�&�	7q�u�Hv�[��;b����A��5ey"���H��5k5�9&��MC�%�G�����G6a�.�/yc�W����p�)HR��śs�@M�ÌN|�s�s���"��rȭ/|<S�K~�Ԡ��KɹeM�Yci>�=��6�"��<�kkF��!�??}!#��fցB��x��Fȁ/�9��a��R_���'����d��E�]���t�V#��om�̇�_\���CX�S������֟ꖅ�ġ{v�p�d��F[R*>W��������C�;��K�ø>6��Ѭ��Z_���C�k����~��ӻ��$����<�:�ЀX�o�}����A,~�������k��
XB�d�j����S�b��yZD����O���Om ����f+y���,�=�SPw|ϯ���io�`����x-���'�q���
�n�ݝ���3xK	#�ݤ�}��T_��8�C��M�XR�ٷv,{��n���N�]64yq��
Qz�B �\�ەHP�ŧ�J@'[�Ӂ3��E��"�n�e���x�FÎ��������[�3;x�RˋpU������S��J
�*
�!狄�m�����a]����P�(F�)p�)�%����b�}l��^6�H~���~���S���bKKT�������g�ff��G4;z�U ��Y��Tϣ�z@�whj�$u˘���薐�7�K���Fɵ9v������w��Ƙ��		���%�z��*���I<�JךcRz �х��j��u���5����T�z�Y�� 3��=le�f
�d%~t�%�q�O��:Wή�,�T�/��?65һ�Jz(�����o�a����#��Y�9�Di��xfX�L&�3�y���,����h�_�f��5�Ŭ]Za��0���}U���s�=�����bQ�d�R��>����V�9ٕ��"��݆*?!������[�������9���͢�b�~OP;�U�x����JhK���AF�(�s��Ӏ#��u����z�����1(S��xAe(�����[��aH�g�U��ܑ�J�}ǃ��{�R�g��4�r�sz��U�f�D3O�S�u��H�|S��1��$u�P�r��T�c�3�<f<.>��g�(p��Z#/��ܺ�G�$�hy��IP��t��
���!_e]��Z/��i&v����KT��_�8��W8�!}�]V; (����m����ѸH�a����{��4��Ǭ�fk)���t#w�����u�xҪ�Vߊ-ᦡ������]����C�H�O���b�%��o�f:s9�:�V��>�pM�}���g�%Ebg5B���?
��<�@���Dǝ�q��q.8�w�]�\�m��`J�>�K���S����,�t��6$�G�04�ذ��=m���T�Y���\F|8sZ(�����2_kh�Q���G�������<!\o��U
�3�^"��km�E�4r����`���^���X�d�!���@����h��yF%d��_�+c�=�ڀ<1h?�`*i��$i��XC
]R���Q��*(?.Xu�q��Hp$eGm�ѭ����H�Ų��^�MچYzz�D��t��2_C�{��'�Z���+nK��6x W.n�?���T������GJ.=����+b3��$M�+�9PO��+���2��.��U���\���DLF}ٲwD���22�K=
�x��]����Z�� ��&e8���O�ı.V���h���$	4�������D����Rξ��3-AQt�w���]�Α���0��b�h�JZ�����>YȫC\>&l����Y�i��e�#�ڌ8ӥ����������f�b<�s�
�z����7Q�u0=����g�ң�����I�tkje��,�a�m��K��K�=R\�2�����ܞ0��}O���'g�L."F�[�v/�Ӟ��SUy��t�S�����b���b�3��*_���.SpY��2�����v�|&� ���m^v
2��w4/=��֦����MQz^߻mJ֐��EG����g�d�������/������&��y�i��Q�U���Xq�<�7V>h:zJv�~���H&͑��dƎ. $��!� ��#οf�σRxC��̽0������@�����"L����G }=}Dn}�>�D+D�y��L��k,�vz�g^Nֵ�h5nVlme���'?�5.�MI.���`����:�#@�0f�Q��c;Kf�4V�#�zT���C�D��|��W��u1���;7K����`�%KZ���*(k!Wwܱ�eϭ�Y��3��5b��V��Ѳh�b(���a�.#e;� ������е�63 �n��E��M< T�IWݫJ+��1+����m��,kbd���8H���S&�e��nDi���`�Vycq.3��1���B%k֯�Gm�}	up�����n�?4��8Q�L�r�f7��Aa�4V�T�89K���V�ǳ��_��o،�`0b=�h�p���� u:<�s�\'�B�jyܩy�@�xr W�xQe���*��5�k����ƞc����S,y�6A�7ʖZa��r�#�w�[,!H��j���78&*�&|0�u�z�{1b+�{F�~-E�e B`����K��'4r���k���2������(]L�!�,;R�J�����?"M
/;�"�)���wܾ���[��7�@�n_5׷�ğ K_ߧ�X�u��A��
�� ���n�qW�R[m���0�-h+d�ΈCE�b�t�5ۤ�@�c.f�hm����D!;)jP�h��^+�W�/�lQ�Z�m�{�9�jjڷ���3B����C`�q���}j�Q 7\�Jis��w�,-�<_�i]�.�	��(	g;�A/��9��Pb��W�if�#�n&�=^�,ҩ�
�[�N��`�38�|��V2]<%2���,�BI�^��O8epK!���WL���մ����g�2}����&&�����^Ѳ�j�~�w�(�!���'H	x�L˗�"ظ�=��T�ʜς��Ǭ���I�	[J/L
�	�8 BL�W�OHa�v_��tDR˽�
ͅ�5��8����+B��F�U��}����{�1J�4 \D��z`w����B���Q��Ֆ�{,��pu�2Hw0/��R�q�r��E�)����)�>�^�3v��7C��%e�N`�t%vx�Bh�B���;��[Ꙕ������f�l�W��w���V�F�[����,��vY��.���]��-�g��]Z��P�����E�n�V+*��js��盜�Ja�?����8�ս
�֦sHĚW�Tإ��&�	���c�G�lA���XԸ�q����e�g%�l���u���v�e��S	�5*��.+��y���C�M�T*�V00h�@����6+�)!��5��7OH�2S�h�G#؊,����
i��� ��z��.G�\G�&��y�,o����0M��ߕD7���!�hx6��3U��t����3��,$��A����y7�7��$�
l.~�tA��;����Q�#�*=ql�.�^�;��SX~�ȿ[�O(�u��S���[Z{�#�V�EO����P۠�.���=D�m��VY�1X lҿ�'@\�X�dmӗ�f�
�,S����^�y��������R�<<���0"&Q�4X���'�&�r���oF�D�HĨ�O�o��;s�4���.6��pח]�#�Q��h�9@� *dO��ה̓^��+ ���L�?�*��Z����Ӊ�]�T�Vhi�+:-��*��:��*ct.u�KN#^C2��d�������nt������O -�W�-bҷ�l�B?��S�!��ȗr-�^ ��.�A���֫��(���~�?s�I�$�ղ>�������^�C��2�O�Ք���=����fYA`���m�:;�pn�"�ؑ;Z\��������ʌ�u���|��'�@��C�.b5Om���j,e�X]�D�;VB<fP��OJN�F�<;Х��g{%�� G���
���Y��k�*�����$H��t�~YD�ݕ�M�,T�Z)sdv�v�90�-m���1�t6��h�Vϳ�*����p7 5���u���Wk�c��md/�yU1.}8 �:���:l�aFϣ筷�ܢ��( ��G��ɻ���5�>���U�.��_I`n�ӧ;
�X����CQ�@���Y�f��^|e�u�7&¦X�3o�pn��6�Q�^9Ꝧ	7:�t��,7��o�����P��Px���:&��D�^��\�4�<��O��'���0���T��3D $1gC��,d�Bg'\�e�_i-��?c	&�g\�Wb�\�o�]7}���q��d���\�P�!͘�P1c�[C�LAHl?����Wk���^,�XJ^R�t�';uC����Wm��I�]�Gm}��N��H���jӆMK�#�A�-+��O �C�Ο�'�yv��v�(�R��p��B�%'��0Y0t��#�e�&Z�,�U�2��/"��nYB����p���M�ʼ�����v�S;�L���Q�0�6��'��Ն��� �M�V�o�~wy�ŕ`���nR�N���~[�(Ν6E�&��Y�P }�3�Y����%l
H�+��&����g�<�����	���֨�S���#�2%Fl��2����pZ��s���}��1SC����l�~���D���T��3% .s�g��,�rv1�I�~G��+�
Z$JR��/C=�.,$���C�j�$�L���>k�{���Y3F�9a�*T�ЉzB�*ѥ�:vd[�mG�|�`�]%�1S�$����QW���pj��Ϋ�ᘰ�=l,^���؝/��mq(�~�ܕ��!Xx�5��ʈ0��ϥ��S�P��FL9������]G�8�G����)�q��9�f%R��:piN��s�/��U�TU���|��"��[G�y�(A֍`,�8I7>U%q��2��d��h?Sd.ׂ	�B�~s���\}�����kO�k�-n��b��,d~)��ce�a�b�E���D���i�R���[�Ϸ���w��0���"�b�PJ�4�R �����1��VyO׍���h�}���A\<��O�?�L�r����=n�=��:��-�Mk�@���O�/��3�H]"h�m��RϹ�ݒ2�(�
�*�����@���5If�� ��~�8��#DA*٘�y2\�FK�y���fߘ��y���]�2��M��1EPD��
�wv�b/$��`�f�V@���U�`B3��?���q4=q0$^�k�!��U�c����Z:�����|��n��ȿ	8B� .�j��B�~hf�^��F�J��,Xt�f���v(SKr5�S��$�Q~!�ӣbŏ&L�e��L���gD�R���g����N]�b�i��=`�ͳ9'jR�)��b؉q�X�Zpb$�`>�੄?�H���K[�9��6��L��s>DN��R͌h2����pn[��,���j�-��	H�'��+_YJ�i�Mo��Y��Nv(��R���]�8q�_���ꁤ�C�Vz��vf�=ڤax-�����F*W[��w��s���r��%4�~K�f��jg�9����}�v:c�ԙ�U��@�P�s��H%��oy�VW;v���N���l���k���aܢ�?M����n5�/�e�с~C4-�#K ��N*5��� &G�c(9H����+(��ȰW! vIM�a�J=hgRZ��e�H*hȂ�S8��iII+���X��졺7U�*�Fy�����g����NRG��!�����j��/05�)�h@�9�DŢ!_!0q����!��S*�j��V�\�vJ�x��D��+�#����u��L�s�.�C�噅j!����Y�m��s������pJ�`7�C��c����+�hBPu@�\=6���|�-���j\4�Φ]cG Lp��'f��{V���i�5�)��;�9��pS~A��n����fi\��3��0�����/�,��Q�P�=<xA��9G{��ՙ/��vsn�;�I~������D�9h���Y�=��:�1u�l�t[��\�����v@r��T�v�Pb�3<�@G�	݈����"�n�d�6���-ż�BW~�z�VJ�2}��Ě��a_6���X��p_�!���Z��J����zG!�j5�ڌ��ہ�T�TH�C����{^`�a!E��
y"��+o��Wh�i=�Wh"s����Ğ���x��6��6�q��,z��J�%!�X�M<q��(������"�60�*��ό�� DV�]���|�I�k@�bڛ	��B�F?�[�6�Q|I�Ӏ]�2Ƥpa��E�y/�y8j�r��E0����jL>�z`��;{�s�f"�>�-�-
���	�\� H��P毂�g��	F��`7>����U�i�-<B��bEli��M4G�?~[�!%u�*4��wS�]�����M��'�P��r��a���ظ����ؐ��������aN@�������V/A��#e�8����\����sro�հ����. �)6	�4��p� �JxȻ��o]V�=�~B�6>+�!��\�3�����wF�dW�umǦ&,���sY�}�֝(N�*T��Z.���(�Z`tP�Ua�wm!3ԹFԡ�?�Q���_��Rd�:�#%g����%a��A&w�?�s�Nk9�tm���t1�X*���������Fe\�et�D��ZW�^�o1�)��H��0�W����&~b��r�2�������d#���q�eՉ}#	��sH�r}�;��H��<š������+D�w5�$SS�_.�Ǖ9X���6�OސՓL�Uq�������{<���y̓����|ȓ	��e+�oK��hŤ���ipi��o)-�|��R������:M&��^D|<E�
6
z�)��.Uk��C1�^=,Z��*C�RS�Td�azY<��H-� � 4�Ԉ�~���H�pk"��c��rOM5C/���
^��+v�̣rk`x���7�k���ϣƟ~ڝ{��	W���Q�;�b#.uA��	3��׋��j�N"��V_����N�Bp&�b�|�0rA���{���>�=��cA��G�!���x�/~6Zl��9�kԆ�2�� �7L���+�^s�t��e�ӄ4��\z	X��@�˴����<�K%�O^ܠ$gT:��_��\b�W���é`�*�ʒ��YE+�m�{r�0�T@�J [�;��q2�M�ΝT�Ȃ��&�}�y�5GH�7�x A���Q#`����I����ؒsb���BeEG��ѱL���u,�a�m����0�Tzw��&�
���+�U�����6�����]Ee|��٤�Y�!I�S��3��	�r|o�vA=5�r@�xx`;�� �����k��oRo�]I��Y���=���?�����Z�Qk�W�F�U(_:�x��~�/Vޔ$h������U� �h��"G��	��ƴ��]�O�SZ��%�m`±�6,R���<�y!U�ă�W�$�����#W!9_ڤ������AQ�$�2��ؘ�[!,z�L$ȧ�����P(��{������d��[86~]�Sem�2�]����}���:�GU�(��Ih�ꦤa��t7�6���RKq��P�î/���ݒ��%-]޺�F1GK�4���z��^�~7��c� ӊ)���ӝ[9�wB��y�� y�#7�믚��*�z����U��7�w})Qo{i��</��>�X��~5��q@�yovW���(�m�K\�|Kcf�z��|w-������w����k��`M�vÔ��A{`��^n�l�T�+Pd{V��v~�ഄ[ˀ�Hi͛|�Ws�͜��ޭ+��si�ѡ�S�L��n�g/�<%+ g�0�!z�Z���|�����ʼi�ef=������u4Sfg��_活=qF8-8�٨��AS7��0Cm�h�y����'O��ӿ\ݳ�|!����4 ߐu4����o�9,�'�fɎ����3��m�!�T�M.yֈ���rc���s��,�t��!W|Fd�q/ōu;�͎��$]1�ʟ�������A{���Sn�������!B�4�&����]'� �^'�Q�|1�����E���y4�3�[-�<�B��j��L�:X�r���� �+ z'صM޲�4.wb�Z�c����"�\B�\�{�h.�G��S�=L�_�{*���e���!8�Aּ+B�)7��D��g�3*ǲ�A۞�g	چ�	3aVk)�{�vB�j�Ϸ�ӑ��h䴹�����0;�[��rZ��0}�?�p�k�e6�݉%��T�1�H�-���L�)XM�O��r�ۘ���,�W2ܧ���N4�:�Y�LeU�����ߥի����7����BC�	�䮄��+c)"�����	���ؐ:t���M	���
��$�Z���gU���w2>%.�k�$�e>�HWNfx�:�MV+_��X�%i�*����a��*����/oIW��
���j%���.��*�'�-�#��W�!����Xo�s<}�M�K~��DWDU�`@Z��P ;Ǎd:<�56�1K�Gy��}��ݜ�U���c@�ɍ�.�g�v�6k����ޙ��%R�)L<�)l����])�>�+da��7*���
b^@�����f���¼X�i&��Ù�;.��,�1���]�6A�]�g��T��](��%��Ŀ@4���x?]���dxZ�y��E�G����}s��(�zi���S��9�v�����^C�����_D�T�U���{���'�{)�V;\����5�P�b6�y$��Hc�e,���t��Ǽß�a�N/�(�6�/��nA�R��ئ�d���Ы����~����"r`�<��'M�!w��yT��L�x�1�=�9(��8<i�����`�F�� ��S-5V���#�nUB�N�t�I�JZG���d��I���,<)���:�m>�j���G�h�Tr-�b��g�	"6x"B�(���\�c�\�9V��-^D��LH�^��v��_�)��AF
b �r���c�f-+��?]9ˬv��~�� 7o�f=7��h�:��m>���F)�Mߡ����B�������.7��HD�
�(�w������񏛢���0�sٺ��������>/&��q�D.��:+C�w���N��þ��������x��U�,N.���z'w%n8�xT��,���'e4�d�Y��UZ�t�4�l�>;�����#o8�&�y����V�Ό��_���U��|� -�3�4S�>|
�*,aq�KrAt��ؑ����'e�o�*��*t�2���dVI�a,&N>
�n��:m��1�?�{�_���[1�J腚���8�e�"�$�@'����^�zbn����^��E�A�E�|���U%�8��s���v!x�b�9)hc��ȷ�k7���Jj�f*�s����a��}�o�9�JM�:�ߧ�&��b?�Q�,�+u��x��՟�j�>��K�~c,B��j�2lvO��`Ķ�{ߥd�gvq�e�
�����_�i��𻬔lv!=���1��Lq�͖�,����l8�7��Ӥ7��OQ�f��$>ӑ�A��3u��� �
;��z"?j�sF���+d,��I�|{=E�i\�IF��H�Yk��E��9ps��\#%[��f�@8�wَy��.��CK3W�,�V"�/��e6�ym��76:;�X�� ;Y�Q��v�Z�c���YW��f��z�5I�ig�8����&�������iKɼN����m"�O�P˳k��C;�V��Ŭ�5+w��"}�Ⳅ���+���O�p\�j�O0����b�>�0���8���Qh���Q�Ҏ<���g9˒��N�}-:��t��1����t!Q�dp���UI�[��u�/aG+���{��)���d5�G��2%F��x��R_+�t��ĉ�H���0��л�K{�ڸ��9V�I�Oۼ5yu�2�����FG�7*����~q8Z��x�~�h3�X� ���%�����kJ��kkMG�U#�$�ޜ�;�&��JUO	��BQ&��P
ڶ���	���`H�J�ggk��O%��C�������8�=Tc
dI"�n�^����/@ e�n¢�8 ��p�|!�Ǿ/��x���r�őa��3_#����M�^y�p���󮤒Y2"�I�@ɴ�HL�,#x��h=�KeX��|�D,a}��W;�~f�j��.��4+���X�ܦmy�Ș���<��Hpx�`�����Rx^����`M����;����1=��7@G1�*��8J}��BˊU쀗� �'{�E���p�����*����H���2g)���FT��A��<�/�\ױ�r����ǟ����Hsp�F���ݔ"�Z&*K��
α'˻"�.����+�3��g���mŨ�z�,_
����DR�����d'�<x��R2ݿ�\�N-i��4���OlRr9mSױ|���j��o�_�������->d�s��O��`�@��`���0�sMBt�W0��K�P�U� ,f�+�TGm@XH~��������9ՒB�B�Ӥ�F�!��FW�p�{ض] 8�����C�jd��l�s��H�4�4��&�ް�>�
�����4�w%�	��)�z0/��^`��yoAfö����x�uϚu,���L���o@��;A�0�ȫ��u�^���u�W]J�gTQ��0՘�ؾNL}��l]��pR�ʃ�/�EP����r�p�QZ�'V}8��P��do	:���"���͘!�|�5�^��J��8�q�����5�i>s�ߕ��O��;��<����{�:[?��b�h�F�ō�H�����33��$ؾ�Oh`�8��o�Dh����n�>��T(x��R�m�_V�v��sNa ��-�ʘ�
�YL��e�����f'���:�������&�W�P�@����:���=-x'^�kC'��-��;J�	}�J�ܗ���<�r�<Ti��(��п8��o�Yz!Y�Q���{��wY�Õ.,^�ŅENh���)dĠ>��?t�M��0:��n����< {oT���'�묒82�0���N|�G˹���$ѻ����^Q�E%�D�Ť��,�f����VG���]~��p|�~�e�$�)��{רڥ��b���v�F��`jA˥� DO\�_�/��w�R���p�O��o�ʞ)�3�>����Dm�H7��:��o�@�k�I&
����Jg�U�m�[|d/\�T���u��R��o�M�ٻ>��.��ߔ���c/�Q𱿟S�����+�a}�9q\����eű�Ub{�v=X���*t!���ٸ��B�O�����`��O�g蹶T�|�o3t�B��׫z��}��apU�ߪ(dY4j�2��:�Ϣ*�<�E"�P��8𘍡2_H�"U��� G,�.�T�H�����}�E����ݑQ^��m�f
���z\8�ޤ��^�(ıem��@z���c,0=Q���ܽo�6���!i�!;��-�(����o%�z�����	n:���eϬ��R�Ү5�ύ$S/�F[�뫍Bݿ�H�ܫ0-��,Uw��&�֋�N8�>O�q�����=�G��ye���n��t����Ѐ��b�رC�$"�����qjST�4�6Sl��qQq�M̦�z>�1�bS��QC(�9]V����R�����7>����<f=�NL���d����C8�(�-�W�rR���]�
u�U�v��&�]h�n�� "
�g�0�Ѯ���'�2Uo�xa������0�"�)2	'\2�����O���JZ� �j��+���k�������қ�s�Y.PB�u�]q[P��C��M��A��L�\��p����q��۾�Kd���h%uH�v��69�W��l�u,�U/VTľJ[��~M���	�xq��K�}���K��{��R>�z}s䴱
�B���S��ԫ���N�	�4�2_�N�l��Z����4Z�r5�::�`jzީ����1d 
��`�di�Z����U�r����BPxq������m�}Ou���M1��y-&�r���+@RJ��v�Z�(t�����G�[�Y�xf����q���1���~������d�Q~���x�rT~�E/�{�ʼ�NGϽ3@�� a��Erc�E)��Ɍ2W��%��������4�&d��UA�IPb��4�����2�AGQ�)��Y[P�;��
Ui-�f/ű�h���v_�>�2^���Ê�xv�[�Q��sWW{#������̚ZV#���V�.X���X#7�5�zH��D���2�]+�(�B��������������Y�ӗn�F����0���I"�� ��gE�d|�%w�����BE"�b�a�����᧑*Lnl��7A��C'�/U�:H��,�W?r��\[����|����;ڟ��)�3���_����5!��ux�M�:�Z���f��%z1�����Eq0�)f姀�7"ue'���WJ?v3�� �k7�(=����D��Ac�w�]��K�?���_hld8
����SK~r[�b�����A�_y#�@�1q��x�_��lp2�!5`�f�H<o	n��YU��4��DQ��S��+5�U�$z ���Ko��޵rE��[/u&�:��}�X���O`5TRߞ|w�^:�x��r�'��x�lst%��R�y;%��ME!=�n�4�Q`T!<�,��E��r	����z��d���o%�wrɪۓN�()��Bk,��j �#x~bԤ��#*����<���C!Z�F08�T��6y�:S�Bzz��vW��-O�\�af~&9���@�-� ��;�tCr�}N3+FHE�|�@�2���h�ԑ���������?){+M��e���4�<�(����MV���-Wj��H�?v�Զ,��F��;���py��7�!�4��͸��I�W�C[R#����������ѡ+�CK�)��<�Foh�*��ebG��xqk ��%�7��A��v"h�����p��c�d��d�s2�=�I09�l�Mԉ n�,�ɫ���ۦ	�X'	�'���s�+<Ut�O�UgQ��u�/���w��=q���ĩ$a�3�Y���ޫ�$ii����m�KX#9�Ԇ�$�/���A�NE����c �b!�Z�b�/�2��I�^S��y�<�J��k��������P�v��|,H>s�y�Y���dsx�9b_��Yȁ蛍����yS/��d?6���.7�\�2�ǵ����&.��*��t*	�K[���v�bC�۸�L>$|2���>jg�z�E�r+Z;۰�S��"yG�&TN��<���ia�uޓ/�����6�6w�r����2���<��K���q���+�M���bi]Pf;c�a-����!���g�&$ď8=�r���"��`B��ph|b2���`�ɪ�m��5@����-�{��-b��Wݥ5@�N2|V���G�_b�鲁H���=�R�ѳ��"�i�^�J:3�s�1��e�8��Br`���w��Y}���"Ԓ@^SoKk7��oV�ͳ�o� ��D�����븪ӿ�#P���T��j��Xs�2f�%�[x~pH���F�^0KU|��	w��9�tx@Z#�$�iI����)�;�}��m�MX��mK�\+�����, *�a���#�>��2�DbcWw$����_Y���x:�ф���,W���{0P�;����	ϸ��'j�BY��E��j-|�1w�j-5�/�'��ϑ�U�-�wӻRX���X^S
Y�"�^�(��B��&ǖ!�C���n� 2``MmU�$~&��ϰ��������t���1[8�w	ɽ/��=��|O�Q��k+�胓�z������V�E��t'�S��Ϗ$��զ
��}����4C�^f�z�@���\.�ʝ8����@�DI�f6)Ci,��w,{���n�S2l����Ud�̎p�@ �ԉ7x����$7++J;��D��Tcp�u�R;�R'ռDM�6��)޴7"�S�:��k}3=Nj���6��X�^��Q}��{�ܥ��c�8R(Ҧ��P���xt���,4i�Ys�|	�0Y<C�<��D���nq�����死F�yG��@e��28Z7�Ɠ;LtKsbe�jQ����� ���m��$閳��4V�_���K��WD��j��/�E��Ay�KAO��F:�2[��+�W����Ƙ�Syf;\f�B��{h�����A駬�{��5f�b��<�xp��E�Z�u�|T��3��:����%<"��d]���Ae&&�11c卵��j�� ��rb�{g�h������ؗµ��+T��ણl�M�e��T�nB��u�>���������-��e��zjޝ�]d�bq��x{'/�x��C�����U�8��jk���u]����˓����=��Ç~�Q�~2"�������׆&�,��������P�c��p�x~`�i�܅w�� rb�J�RB�'����_��9���� eL�'���Ec��M9!��$C����n\6��ҰO��Zi���lY��̴(�E��j}��rӴ5�]]�c���� �!�Zu��0��4�@*�Z�P�p�U#��h��ސLyZ��1��:C����ka����D1�"�䡇��n,�]6� W�JQ*Zi��{v�r0�Hrm�4bԸdi���HK��XDdZ@�?�i�Q��.������/	���VO�_x�'q�=�WB��7����U���'|�k���X���He�����Ӓ���E�B�6*�1�+%F��ޤ�/�$�{�;R�����8I�¡DN#S�,�:,W�T�X��n�.�`E�8��㆒f��N7�d-xb�H�Q����d���#��U��;0	�w�O���`
��_��L��yE͕֕>;���O{��F��<�Ԓk`w�7'DWi��t*&��)-�U�G<X���wjȶ]��^]ʣhlB@E1�}���3��U�����!ܚj3��R���X�:�uO�ʌP}������Pd,�Q�#Y����{�����7?$������#W�8@�|�1P�^�s6�䊷�cם�p��J��K�Ɨ�����<�iם�ᆼ�/���?���.��)�"���� �����.e�ލ���>v�H�b$�>4����0¼�}�Ch����&ℚ��\d�v,��L�׳b���) �V�Hˈ7����1�D�f��i9#���\�B��_���սm���aĩx�4�4B��:���2��<O~ѻ�c����d ��n*�*m�5�Fn��[�o4��!X��~���`����,��褙X�
��3�mn���(�t���\̫Rc�"�P�c�u��vy.���1�5�"@�|[�j�k��Ĳ�	0�v"?lmr�0cs�����W�"r������;w�A0���6z��
�p�lִ�z)�\q��,8���_C͜�hD;��eE	G7R�WW6/0��U1�(��U��ɧ"fm5G�*������,C@} �?&�$�%<�o/�EKu���|�#�Ē�sEO�p.��h�\�f&��&�kv�A���n~��g��>�v��ˉ�\��^���2��p��_�^���n,���$��=�i	�0�W����%~"\�h�1��Lm�	u�^��h3~�����=�@D����݊Qg��t�q�2dt�`��f��$�ɒ��[���,��D�Jy��V@�����`�T����K]��QIϮ�w�(,���B�C�-��@�$��!�'P��;�iR�8��PD}h)�U] ������U6Y�l��[=KFT����kq���N�������|�[P��ɵmWߨPf`��T<'�%�ͮ��Ĝ
)�c���<TBѲ�IPMh;��QN�N9O���i8Dt��p��dW"S����#��-�k��zY ԘN{#�����g����ʾH�X���+6��&�8J���H�3*�h�i8I�X^��t�M�Xб|h{%ȃ<C�'Fí�.+,���I�x&ànZ�^>v�L��y_�y(&��}E��׎�#��I7\d7�x#�c����V�W�U���L�k��M=N��I�A���5Erk�`{��F���a�U	_}tCFRV�}�1F{֦h�}�Զ"�|=ۙH� �$��A�|���~�׆�O��p+@���pH(���������u7�O���t��B�_�SAn��2�����Gx=KJ�u��Zl���
�J��B�_V��\a�џ����b�Q�s<;1�񄶰���T7�:�ׁ���-�S*ϱ��{C�JV�Opm�
�݇3[�p�tA�O�Oj�*����4W���ΡB9�Tg�NTI��w������
�)<p�Y��}�u��_�"CJ�V�"�f�TwB��D�C_Y�(z�[f��F�����#x}��}0���޷�k\��P�)���R�5�WP!�.X��y���>;�~!w��� @|0�S�'��j�����D�ATD1�v'NBƬ��B�l���M������U$
������x���aQ��	�#ə�L(G��|)�a��j��$�l)���� ��L�φ�~��1��i�!��M�x�v2�9��y����p�˗�SR��x ��hl�"����Î9Ŝ!`qZ�vչ�<e7/���5Ʃ��02�h�>:rP���u��������U��o2>�e��rR�%���V+<В��!����{��[b�²Ғ+�9  �����A�vJ�冎��C�������z�ښ�� Ф`�}��r����� ��A:�����U]0;Ȅ�Q��ܯ��K�t�1�%������R+ak�����r^B��2q����t a�^��了��N��eYk�0�̈́�-��ײwE2�$�X���Nz�Q�FJÏ����:G�a~��æ阹��>�������XJ�����u�C�
�n�=��~߬$|�o��� ����mÃ(�!卒���qفҙ�cWQ�:m>� �a���f��_9(yF��ު<~~�0D0�5�X�V�1�f�%3�	\%]�5�� ��K��P[�dvEw�qU�:��8\Н+��ZYu�e���!b&����'�"�Z2��=Ҷj�eZ����<�\��
q�Y������`�x;qR^^�G�q^j<ž1 ��݃H`<ؑQ��y�a�Uc�+��U�����Gu��BA�)���|���>���01��
�-�b��d�<�&$��Ws����Z��w�s��d>�����*�_�y���O!��οU��h���<��l�n��������<�#�J"^�V��OY���&x��r�1%˱��*�t��P+�K�h��P���c	��ѻZ�=��k��}�n`���ܝ��{@O+��
JP�f� �|���r���PQVg��`���.���7,MR���^U�&�ٻ|�s�2@�6ס�~�u�;A���;i��g9���~Ч������:!cÝ�k'�z��Ƽ�1���^K�8�;��Z+��z�lC)?$U7���Y��e�7�~ ��n�͢��3���7vk�8��y�AS`a[�����Րu�����d#uܛb��U�j��e���,��E9��u�}hĚ��)�|���Xք��e �$j�c�0-o��e��yǲ�?��N9����>�����$����C_.��m��Hz����l���
^�#��7}(#�����@�$�8��A\0l���gVs&��!Ic�ӭ��<�*f�Z�d�g��4��߸���������4XR��� r	kׂ)-t���@6�So�V�D��b}��UW�%�0eѬ�}rK�<���Ii���[%�X����1{6#+��w:[����Y^�Pn�n焞`�9�� �9 �V�ޔ��S����RD�Dy4�d�n��\H�P��ܑ�i�*���C
��q�_�Տ1x\0�4���Lg~��
3x���n�p��H��ÅJ���|c�a
~0Zm6�f�Wđ4�n�"#k|`��o�<�_�i��ϖ���b;�~r�=�����U���%̝��|�E9xa��!���&�(.ze_ j�v��K�*�'wX�f����/+2�&���2Q�Fʵ���@x�J�����d_ڄ����ߡ:5s?��2�G"�6�i�$1K��Ft���Z�2�k�Ś���
��>��4 �����\�^��L��2S���E�Mw�2���*���K���K���AKLRj�(՝嗈l�DX��4��R�/vx-�*��㩒��3���s�O�O��{�C�b�#ܙ��`�a�T��]�KvŊY���K��6��AQwL��3�s_
�J�6<�U��%�=
��}=�e>�J2*�1~��p�P��M��!���"�+;�T��������!8�{��9e6�kHF�5 �5�B�_���a�������Ffv�rFP��k
��^�t@�7�tn���A�p�-�~��Ho�· ��s�+�\�,S��l�|�`w�)�<mQ�<|e� վ�4�U�'�ɤo�/^͠��Z+����X�w� ����Z��]�jit��$[�0K&C��ɸ!h�<�\�`y�oyk^ʣ������NB��E�ޣ���	&�b �[�G���V+ˡ{����� @�ÿ�܉����T��v�'���b:�k)��(~s:�#R��腮ߏ�l����W���%��K�G�3��:L`y��1�X��mY�g�u/x�r�����-���1�*#����D'�=B�,���!�_���԰��]� ��{�#�L@NͰV��4U�����mq�[z�d�����?�Qp�wS��"�&�J7C�7�sz�<ê��!v:g���=�m���>�������"����<0��.5|��\�{��m�n(��ͨ��lIL�T��S"s^���+(��`�AiF��ktz����Skg��ƴ��.ӭopX��J4s2���B�@[���R�Bq�����Y;�P��7l�n�{��-H��-�TC�U	�RI���]0S����6!��)��|J�K�G|��gl	:{W65���}�ŷ(s:�:Q�1,��ꋧE��rʌ�D��@=A/�����t�5&�n��)�1�9��-��6�3�h=�8�WHgG�h!�pz�	�L��=@���� m�p�o*�|M������=.b��U֢U�aj:$3���5%�AI�0&�`�эiy��˄��M�F-ד�s����A�!� ��:��߶].\��(�fF��w�':������`qE���#�b�@��D��gI�}��J:��F����A�eƃ1W�R����J�8�2�������p[8"�r�"P�{����h�S�ou�,LV�6�)g�u�i51�
�+�c"(���SƃG�{G�ߒ;���ɇ�1�M���;3��i�j�S'����9>���&p��$�Br
>��.��y8��N2�z���S]+j����F��%AD�V�Ŵ'�������VQ�{r�.z8T�=m��S�����DΞ`���Ij�eJ3o��4��pltu�>Y�5���0�ߑ��<��/ ��,�Azz���<��qj�U' q�Dz�����"D 1#����䔷���?zU��afo��A;{�p7	�nJ��������iNc�~�3QAڰ>�����Z�{ 6�6�\C����юL�y�h�4E@cy�|�eI� h�X���b��
�bK�=G��f͟�P ZYczg���ۦ��g���ݨ��n� 1n�M�'�c�3GR��*p衿_��G-�ex��$�����z��8&�k��=H�pg?�\�/՘8K��ݦ�
��vD-=����5 �Ayޑ6�Y�`Ȣ�+��Y�C�p:����6tV�0�	�ǉq�:�z��,�U���T�b�#�G~ҤT5;B`�.�WG$uۄ�0��٘g�Y�l�m������-hb�:C���(�)rhm:*�9�<������y2���B/OC������s�ZOoR�+w7=N5��%�� ������&�L��I�
u�7��xm+�Ib�+�S*y��}
($Nn�xI0C���ﶻR��(�*G	'�Djy�&
jۼn�[eLiU�ʜ6�3�D��b<�^�]�6s�L��y�%�B���/��D��|�V�/	�r�����eGz�v{崝�?�>��zOlԛ:��.���L���)V;I��/8l)�!_��5o${��xEՈP��r:8�(&�0�1 ��H���2�4R0�B�1������c��%���˩��Xi) v��~iU9B�	}��6χ�买�{�y�z1b���w'��#А[��&T����F��K���>U�����Ì�f�t��p�;�ÏKK0�����+_��f gx�s�\���Յ��y�d7�%�����R�XvŌE��~D�YVhև42�P�e=o�w�12!P!�]�㓇��o]�H��{T�&����%c�l�@�5}V�����:�E�q,�J��լ�_�k,"��x<�f�g�B��P9����\���� ��\w��k?�*���ʻ��H�S�Ţ����j�2?��l��$��G��אq�t��Qc�uD嘳�7#L�p�B���xv
߆K�(�U:�d}���@�Q�$�3�m� ��ͩvVDaĽ�s�v��v�8�_�C�u�Y��ev����Y�d1�4��Ϟ@A��u�B�pQA��+��r�h�Lƌ�eq}�8c���P���twϼD�`LQ�)бw����9M��#nd4���:���D�_��$�EfDS�>G3����Dܧ:�5g9��	y��;�0�2?0.CK#?�솃��>�v��$~||�����\�!<�\�6� ڷ�r���� �8�y�ʊs\Q_3�i��m<I��?�	�;GO�^��pT� ilV��Y)�ږ�*�j�s�����Z��D�(�9�^?�gk�u�Ջ%~��liˣF�u���3���.m�F�c� B��;n�ViR��Sf�K���-;rj�!��:blywp�,��l��-�-m��ik�kH���0����Ѓ^�^!儿���T�/^�a'�y$�p�ǆ&������z�JH�~Fy���N�&5�N2�r:������l�	l����@hKDOvI����`	XDM��Ô 
:��;��J>��T���$���x2L�i
�k܄u��@��E H�Xi���U����u����"�T�>�脮Tj�H�p9��1���T�h��o��0��19�%$y�Z��*�ɱ����?��6��s?�eH7=uR
�7�x�f�)ɬd��s ���A�)���r]V(Gx]=;�^�����&#J^�[��� 5~��&�(����XHȚ�3�^60v��'�0��:΄{ͳXܧ|�o`O�A��5A-ܯ�z;�8���P@q�p/gi���)��<�jZQ-����(��@�§XM�0��n~��hE��p�{]����97VB\O������#��ӅJ0�fa�d}��n�p�������vspy��:$"�s�����y��L��`j)yZ(I�	�O�X�b�&1t��O]��2I^�V�7~Q��U,�N�L�@@��*gp,"�ב���9-�'Z@�T2C�*����s���)6'�i���fy�����C��2D�i���c�U�׋��D���K>6��<�5xKN�����3��r��O�T����y�ǖ6<���є�dA ��9bKqo�a�&\��ݣr8�M��:��	<B�ʝ<�Fڍ&�96�,�['E�C��0��ǼS��R���/�٥F���>D�rSI����a��k箥�:���U7A���P��տm��HxżL8�R؜"�FG�a6��ȫRN�GVW9�N6}��ȕK�	�E���*'7aA�78<��=���N�B��i:� g/��9y�l�Ҧ����� �*����do���$�	�9���^�)�IEU��qB��M�V�"��Vݶ�a�zC<����a���t��.v�['���e�t��=�o0N�l��	5`^2��/�;Xykv�y��3l-��\6��
�|N������Nɟ��K�>�#���t��y�֟��2��*���T��so���b���IeS
`�6(���l%��._�O,�X��f9��: ���vqh�I��L�ƚ^S#�\+�w'�m$���9�>
r0u{_�����_�f�lZ��Wu*���~@^�x���$-�?*2AU8w�{��pZ���B��;j��I8���7�LrE� �n	k~Z�#cN)h���m�`^,�>j~ ��_��.��<0 x�Hm�_l�c��th�A���	���G���
�([v�8����iJa8���AQ(ۄMQ�}���lZ�C	��sp�S\�8�^�Ŕ�;E��������j�#qH��]�=(V6@Ѫ���k�CJܨ��[<Tt�*�(�[�ʄj��K�����wM�<D�u�N�z5��4I�JW���� !a������k����L�M��L[�K�M5���w)�Z��$WF��	��Ӕ!�*ęK,�j�A�A�=��8�MκIө��3V�����*����1��Q�!�-g�x��u5ԆB���9/+m7j�}��vA�3D�9�7x��6��L��|�(
����-�a�rr%��EkW�xGr^�~ �>96sίf"C��Ol�8`7Z*�����:�'����#R�`؄~J��8�\\���1��+Vɖ� ��ǯuU�%�jk��	�}�(��u�7q�]��c4�ׄ��f�
 ���2\��},}�_���8I�א��䤤��C�m��-3�p7u��O��1�uL*`]���������#�yJ/�*�
{Ρ�%V�k �G�U~s�����9��]�l�z��e{]�����	A��xU� �\"�;H��	"�� ӣ�4�`B��`�>�t3������0h�����8ѣ�Fojˢ�s5� ��@��V�-S���xfd������-Ȃ)��^Y�~���|�ؗ�޷`��d?���`�ѢgP�
�8�ӊ0���\���f��߈�Ʀ��;'n�OTjk��ƙS�K��m\���2n�F��g��]�Sl�����x�s�B��y{�3j� �rqQ���e,�~� �C'�sp��eeH37�=�k��D�ޥ���>WݖSa�����).��?F����dE��o�}��{?Û���|JӸs�Pt+.��m[��&f���h^Df���1C��������j�df����.P��b=X������[?�G�5����n���^�'���Bl�
���H#���(�%hύe j�G�'E�j�m����Aal{�ߧ}�0��>j�{�{0��#Uy$6�{�%eP7
�*�qܐ{��\�c�eԣ���O���	�pz;���|��iQ��t����⽄���k�q��@$㐡�Q$�(�/���"Ұ\~����8� z�`�ϯ�����B��;4/�i�q���P"
}O���:�" B
�����nE}HE��Fl�@��r1��QGl��v��gŔPi��,X̑�ی�4 ��4^7p�X�5�N��p�(J�O��5.�&`N�u4]��[��$o.]��&ƹ6 �0a?Μ�^G�WR?���.7hɸ�;[ R��ݘ�
�����}�3��YB�B�N��+G��� ���T��F,a�j:9L�M^-��s9���'�K �b����Z��M�SASj��Э�M֡ 7���S\��b��5?x�K<���+��ټ�I��̆�v)�aA,�L�����y����ԇ�������$���w�0w��VA�+V.~դy�BH�h�5C�����5O���^b�9�aM{)w?EaP����D�2m4I���(R��?�{��G��Y��4ZH<�9���$v��(4�Mh��<��=V\Jd9�&� ��>VT�����tN>��n�7�^�X^��P�n�
��4~�B\u0��!�"5e��jT�r��ɸ >\Di�Q�|b�ku���{��}�=\H�pf��M���f��y��	���dV_��؁~ヾ���r��y���D��G	q�ΧHǋ���J���gZ H�82�:M��Bd�~��������n��?R���z,Q�'���D�d�e�^��vn�ם]��8�i~�� ���k��.)�zs�G��*���2�c�O��Rc��6/A�C�\���fI�5Y�oTCi� �}�-�>�`������D�]�{f&`����|k��\���x��+@B�ė�5W�Z��&׉a���ٿδ��@6NG����Ŏ�d������J@7��4�°b�)� |d.��)�Ge:i�J/�0��;�Z���I����?���\Eǵ��SY�#�*��pQ$����>I�G�4���E�V.�~�>�nQN˱a�R������K����'�Is�o�^���[:akJ����=U�q�?���1,O�5��$>�W����ح\�#��LTAcZ]	�d�6��I��E���xR줸W+rT��/1�q&�O���Ұ��۱C�$��/W��yeC�8x�k�*�Z0FHi����.5bJi�:6�$�o%ܳJ�MEY��}��	S[ӹ@�멨s?��'h<���
�b�u��蘃ӹ6�����pI}�p��p��u F8���4`�h�Ru2XL92� f6��Jb�VC����El�s��Cn]��:���:��3��i[�It�g�r��q�/�ˁý�A�B~}8�"y�h�fgT���;�-u�x"����V���H*s+�ϝ�r�m��{��:�����=D�ê.].��,v�E"�~C����6�4�K�݇����������4yT��U7��6��uc��ad���J���d<>�H�&�UU����ka2��°��1Wh�j��E�2%d��>�0K�֞��]���@@_�4�Ds�v�V��Q��`ǂ:��B���L;�_ߖ������s5ުe�?@��t��$a�:�S�4��F�J���G��﫦�Į����q}W6�xf �!E��F�"3@ 0�.��tF���T��F��׋C�y~���)�Я����AosmC�y^�#���7L�&W~��p������\'ܱ��/1r��U��ȷ>��H-��[���[K��֫��_66C�-��+qp�H]��B����p��Iг�(�6�nB@����0iK�ϼK���;X׺M�ɪ~���OCK6���FUr33Ӗ��V��%� ���ucZ��M῿��W'�zY�c������9�������9��1L52E��E�.8�T�s׊���g��7r3����כ���XA�����	kQ�۵+��nQ��
45q6�%t�\'?�o��3��n��fl8�8x?���i�h���ǻ����.0Ҵ����Q�k�T��|�s�I������W��H�1��ٱiang��w�ޏ�T~o���z��a�~�;��'�f~֩���zku	��7 @��Z�<��{mp-]���������{=_����AcgԖ���W�z��&Kg�S�=.��I�A��m}2�Vpy6��ٰZ�Κۧ�t?�k�Z50��g��2դf&��_�����!�kI֔w�t3(j��φ��,�y�N�3޵P.��=�A�����+��ήRJ���~:��Zm03��;�C;ߑ���8�l����T�Uń�4>,��K^! �Rގu�?���|�r%�bc�yh{�LB����t=�WF�U���:�.�:���#~/�jYP&��OJ��=��v���n[�M�>2N���"zGbyT��	b�E�[Dwb{jH���d�h:�g�7����y������q��]"3�N�|�t��xpf|������;�#�<�g���V�ʙ)� ��SV�"� ��^�����Xt<�Cԁl�Ȥ�6C|��Dۨ��8�p$[9�Bn�@���?duK�M�o��'Gʨ"=��>�\X�YGB.D���u�^��:�b@�H7�0�	�~F�qo桗��T���mCAs:8:�2O{�����0�G�mԮ\����9����O~��4`m�S8��gT��\E���=g�>�>;�k��<�	��َ�����ň\	��y�bv%� �j�M�B)����n����my������&G'��(}w�0؈�Xa�u�&�aZ|��7�n�hf���t~Gq��^��RCub0�WqD�ْ(�.��V�۳|����d����(ۤ��pKV�zq��MN�(���H����R���}`�J�+�2��C���dSݖ�������e�	QX�%Kg�'k2K�#�{���lV�]�!�ph��Ҽ�<�&FxC��$s�~�3�D�ͩ5��,:�5���:C@�7af�8 ����9����{	�땬=j��k�&=�q�Y�A�|�HD��뿲v�8�����߯�G4H9���~�Y�>t}�c{�rb�ظ����g���5w����W.P?:>�m���m���s� V���S�R�W\����w���<����?�>��	�;E�ٺYz�3��D�8$�ScX,�\>؜�m�*���H	)X�C/����6cʱ%�|s�d��R�҆��=�틒��¾�L~��imk��Z�����m�T�"_s�Q"� g/ڟnI����
m|����^��^��	���%:U�$0�
�0L�{���Y@��oOu�h�|�,�������+3��p��"`�Z���p��l-h���ƻ�ִ��?��?$p�.Ce���hf�s(7���xwhX48bi4��=N_��9��އ�?������<�/2��w�ĪP�ۉ�qV��<Ӫ����G��IP2;f�#q���묶�u3O,'־kv��a�� ��S�TX�ܥ�pi��*�ӟ������������RM���L�B� �e��wH�h|4Cc��u�=�tς�I��塌�]���c�6{�|h/����Zw�����Ĥ<�ʝ�4���tƺ��p����q{��E�](�-V�9iM�]���1���������G�:j���d.�H�.^�g)�fY4�f�M;�%'�𴌊�2�����Ԝ����ˉ�e`���u�'��n�c�}��YNXA&��I?�������NQb�x��/�07�}�D
"w�z�,�	����lQ&��L�J>���/�GU�P@lp�Xz���(LCO���>C���Ke���g~D���}8�h�x�/=V8 ����aǏ4(�P3�[��L�A�f7r����,O�m8�	������^~�y�xI�(�z��h�oU���e.���r��*���T/92�[��']�r�� ��ia9�{@l�XM����ߑ6 �rߘ���9L�w�l;-��'8�"�^� ʥO�������9\oed����o���[�B� e��=�7y���uV=ˤ�Z�X3D�`�꛿_�l-`F&�^)l��j����fT��'ÅH��]��ij�>���f
K	9�UG%Ľ�E��L����r{�I�hc�.�o���)}�1`���+������K�mk�q}u\CS��$k�e��R�)v2
yJ��kJ��S���`�۠������(��T����� Kd����'���# X<�X��F�P�@�����#�/N�U�v\���r��w�S�x�WЍ�	��W��(7��_{�T)�Q��b�$�}fph�Z�N���xQ�yg�V�Fc;MU��t��4h�x��󖊟�$)x��'�K�,c�-�?�9���ޟ����x�2[W;�%W�ov����m�#��E���
�����F۸��z3
!֒B��Qn�c�v<�|�1c�a����O�(�=� S��L�q��#5��)�W>�h��$�ᷚ,�	l��76�f�R���ƇJ�����������?���Y�D�x�5>�����$��~��T�n@����g��͘�)�Wf�U��NT���Ns9h`O�@��<��:z�jx�|H�?�U�����i�����SUB�
��6����C�����ign�?>��#"��ֻ�����'[���΢��]=t禝.O!x��Y�\]�6�����I��4�X����8�B fU�bn��gO���i�Z:�<��Y,�/�e�֐|�ʛ ��w�}����d������׎�q�5L��Z�ӳP{2BrH<��[n�ÏG��}b�r�	�P�S0�	�,d���c�ީ����=+����ɣV����0���M|_�j�cdMg\��b�c�b#PFo7��Ad��RjM-Q��,���Cye�~F	��{H|]� ̆�F�x���H��L�H{{Y/����Z���d�]�&hA��2��K�̦�L����>Ns�kB�J
�/�=NM"׋Q
�U�����4BZ��DP�qT��+��g�+�⯕$e�F�7�ւɸd��b��i�eb��w��~�Dl���t	�3�GZ�L[Ui�tն�)N�^�J���~
�-��Z4j)pf�&�`��BtS��5��M7��qx�̲��=�w
N/m���Zv��l�r��9�|��*���t�Tb�f0�J��BpԴ�'E(3����}۲����SѾ��G���c��:]����I�������̢F�w�5��~�z�ə�J&�dp#�b�b�"%�[�Ǆpn*pk�=_�'Y0��3����|�U��� 7i�W?��}e$qq�BЮo)�)CKB/���bi
�y�����?�R��a���Qu�h���a'M����KzʈV�9��;,�B�햢o�X8�ds�ɵ �ȗ�ظ�,�V���t���7�r����*%�]�1NT�+��>j�xV2p����ءQ;?����=X������r��B��|��|�%���=��`9�w/��|cq�XUN��LĜ },{��?�B���gX1҄���s���NgYe3D�q���^�����WK��=�=8}���|D��A�����R�Ӂ

��[�`tm���cEd��"aJ.�k����0�*oX�=�Pg[#)_D�N���L���$Fx3�A�s{��LҮ!��8�oq=A����E[��j�Ɵ��6,�x���J<@
�wѽ��$��0��w?�Zx��٥w����rx�X���^Y���ͧ&���"3@j/t"N�~��"�>
�M4�u���Lx�+���U��jъ�R��np��F �YT�U�����)S�Y^|����=�x-�;��Я�z��ޘ1"C�z�1�q�#΄i�� �pf-&N�}�`FE$WZ�O|�z�����AEx�Q�L�z-�La��93�7�]h����9�<��Ih����b���\���J�'������ѱ�*r����}#4�6~�<�_>�`���]� ��r��.L��7�!���4QH�4��Ua��8��m�E�<a&6̩\+odw�}%�e/D�<��Ǟj<t3�@����2��V�B�@�����3f��܊��r�=�w�X�� ��d�?�q}����qZ.����W�=O�����j`'�qӅ�}��K�6�л��PM垘�#$���,^νr��H �-����(�̶��a�3zRL��ȕ&���5��^��,@� %���}#�ؓ�%�Ӵƥ@F��=��p]DdaÚ_�7W}�xu�_⳹��T'w��\-}�u���im���i�g�T���@P
1�m�9�Z�Q0e�Yq��%ì�J�'[PE����<2&׈֪�����ecvE�N�6O��i�-����T!%r���U��b�pyc�|��=��a�s�a�x�-8Oi�%@c��[��{��������o��Z��"��k3�E��w��2r����N��r>�.Ӳ3���,�"aDt�aÖ�r��=��&+��Q�v�&%�;S�Y�[(&:��8"\J�p�r2=e�[=��R���H�������+ME$�x������tr�n�c��,&/�)g��R���|P�����hO_��~?�ث��%��Z���=B��ڥ�1�q߳����9�{�"�	_�ڣ��T�#�Ac-��_�U�Z�/����aػ�A�Ӯ�[��`��Ђk�$�Y��`,�/��+Y�r\q="�J�]M�P�M��M���Nc�&�$ܣ�����d�g�.;�M�����B����dJu ϵ'�^�%o�ݼ�IW���xXyO�!�G$������e8�lT-�	�ʀN/m��ڙ�H�V[N��*t�8���gFs ��(��xȦ+K�d�[�Vnh�.Ao���y��ş"6�*��Wi�#tH��z�
�u��l݉]y�<�ގ����`�k=�W�����>3G����2�x�9�]|�
PN�Q�W�t��2~?���"� ��~�_G6t����=̽�Z��D��#f�O�%\�w't}_/���;v�/�g�S�HW�ݏK���a5?Y���`��n�o�Z`7�b�
�W�
�\@� R��k�,��v>ժUk�>>���x�`i+��5��ECi5��XǊ�\ JT}�-���~�&}�s�3�H7��é���ǳ0[����nSI,�;�dHw�≾�n�*���� ��Qh�����+�Ci�_�'��lCUc�s��J&HtA,$��2�ڐ��z�*BD��F���ˀI��{d�ġ��e:Ͷ���n��3�	^����G)mF���QۼX��]W��b1�MJ"1d���]c"�Ғ <�J� ��]qq�3�9���$��P�3��n��A�%��E�U�	>V��$SyZ4���"v�n��\'�40В��.���om:��a�j�F���E"���sӃ7K��7��^�)�@�OlL\�gT�%��Y̶�N� �����A:M�ͬ�I�l���~�`�׆z����J}n���'�f�c`�ۢ��H3;P�T�	���ØI����,�;infq���4O�Q���������}\��!�tƚ��d&	LyҖ0�G�W�p���B��W�('�3u$���2�1t���j0���]�C��9<�:�'�?�e.����1��N��?@�f�4���=K")2XL���m�59Ӆ!������#%i��AD�2�#��^��/�[��%��B���Hw�:�yY��q�b���'�9_gHJ��a���o�T�i�`80��.��&W�$���i\���R��Ԯ@7�y2��� �f`EV����7��W�BZ3�(-a��4�US(y����=��`T�]�ܘX>�)�w���ްv��G�F��������!�����C��@�nA�ӧ?~�ҍR��ڗ�1=d�{[L*Ja{�΋~�q�CDR暣m����*�����d�\�]X�1��AV�x��'8��S�Y?
����F^C�h(��8�w��;.��
lt�x����I[8�u���܄�t\z�[hă>^p$8rR������.�x�V5��	>�;<{�B�I!6��0�z)�����]�x6�Q3�1K Y��)J�YN�ۄ�:�������?'P��<3f؄m�4,�R���JӲd�[G��HR-r��d#�����msE��b?�Gl�g��s���G�p�o���(��?�yK� ����l�F;b��毜��PR�`D���S�@ ?%�F�g%�G�w�
N|�4P� ��U�Qh �}ې��L��_��6F����u��=�@�b�� �CJA={Ճ<��2��Y����WO����s^���L^��D	����iap%,_7_��m0��Y)M�~q���y��	�2@p�_�^�+�"9"k�W�&��^X��<otJ���G(_��ϑvG���΄�E��=4!�+Hl�r�^��]lc*Q^=s��b�ɩ
 ���w8y+�/,EDP��@#}a���J�,�B�\�~x�n&�0&�W��'4��"�ppG�ylQ�vE(���',��]�����r�!�K�I�<�a�J�$��_Q�p[�)DQsi�-$!u��	l�l\�2�q{GJ�~�	�7�r�Ѝ���iqp;���(�ͻW�>$�9u
�o�-�E�C@��L�K�L׮Mǵ0��^m�v�F\�F�<|Ob�Z��AK4��9�퇖L�юH���B�`66���`�oK�}����PM�7I;4��(#Y�'�7#E�������K���Cc�\�Ge��鎯Վ��f�)�(�w\W���p�!��o�Y_�	0>�R(�$Df�f�]J݃b�AˡM�4E��0���Q�0[Lz,��@�=�C�]su`��v���}��_M�|F 	4�-�ޒ�z�����3�n�ɴD��Sqj�1$v�_D���z�\�P�%�DhY�f�DJ�ʬ̸ ��.z ����V�iNE_MB��v���y���Q)��&d�v�h�����<�,������^Z+�a�X@:x�8�O����J����u�/�&0®邖��$=�3�9&������W���%�euE�	eLi<m�f��A
8i�eZ%$J;Bpj��R�o�&Y$�3$_T4b5��߷j�E ����Y��	QW��J�X�N_��[�D�Qr�h�ě�賠���|Xy�鿶���N�ͧs�rq�V/ER@7E��ik��殮O荽#�=�����cH+f�b����?��>p�Q���b�4�$�z
��e�4*=���D�����к�݊�}�����T��s�(��L�����k����^��	�l��_��z�$���h�k�9�9`�۴ �������pB�2%Ó��ȠO�k��=�4�`�{�ʻ��F&��0��Z�'_�$~���(�A���Q���A ��3��lu�i�>!�������7eAn�5�����N��iP3�O�S�
�JP�kNM���G��=�KX`2���|�G�x�������4��|aL�������tx-tyY��noD����ωI�g��0����('��UkYK�<K0�W�jw��O��ӗ�W7}x&9s�}��zۢ���"�S"��[��(aiĸ��_
�R�����&Ym�KV"q3�2%֧l�NF�\lN��lʛ��Z�*����q��	W�N�6��Z/����.(����xj��h�J�}�ҕjiHwC���+K��XӸ�䷀zNꐫ�'T��{O��`��et��aA�P���1�"xrk��*a(��0j@4�.��2�"��s4xO��0��ȬLqMG-��K��~�<
aI�y�r��C�$�W�[k��)����Nn��G�K��J(�`L��y�+�-?����̣�K�����u<;T�鿦&,{袝����i���J�_!�hY&�W���s��' GT�߶RA�3��'��A���2�υ�Ԧ�#��3����`-��ޚ>[f�e���c ��<�T�k>�ib�h���q��1'�l�6�M�7�n�2���)��"�&|MՐ�j�W��}�`J�3^"|�;�	�3�)��ɛt�A�$D���ѩ�׳���{"@a� }(��"J���}�_���R��f���gh�y��0tj!ML��=&s�U�a��F�+����z�5y&�3	:�,�k�[��{R�$�F�RN����>�(��;�������t�z[�r��E�H��Ye��@�~G,��~�y��ɝ�B), r��OP�=]'�L��J�n[��C�޺�nv����t,���ĭ<m���찗��ո��W%�w���<\�����?����X����-T��:������U�+$71yKK)�S#?��I��ԍsYdpUD�l��=lG����<���C���,�%���,�a���,N��s��0i��i��I�܊y�A��HH<�s"De�uUK��`f�����Pԩו_������v��=&�9�Z�m�_??_�-���\p�4��S	7�WJ x�ùf�+����1�A��Jè"�%��ϐ�;�Z�X׉I7*M6�Nqj�~�����\�����R���$U]�H����zF9Ďۄ
�&���dZ; �yXXG������a�dT(��o)�< ���@�A�U��p9���;.���OZx˂)F(�WI����o|s��Ah�(��i��Xn����D#���5� �3��g�q��V��f$�x	��F�c	KR��8!��ir2�Fq�Y5��Cp- ���'�����v�&5b	���Fk�vp؎{?2������b�Њ��ova��~D%&�\3�̀c��7�������x��b�o���j�2X~�7�_�j�`�I�S�^밠)�`=��kFn�Z�	c��*�K��2P�n����+~�z>���p��b�|����6��4�� >��d�]�S�n�6��]�iS'�����m��p��J�#�t���p�ڿ��y�N��0��_��sC���,D�����������f�뚃n�V~f���i���~��� 얕P�p%��Z��2��e�1���^���D�3h���=яJ��8{���������9W"E�0\J\Q���20Q���._��C��k9[j�|��A��]&7IP��Ϸ]��r���/���B"�$f���4~J� �q��'��rmm��_x�7c=�x��H{E���[���Cm�*��dZ�К�:�ָv��l+�� ws����1F1���W��>�QA��+V�d+���EYZo�	Ⱦ_q9�u�5�܁	I��{���.�I��H�A*�/E�������O�݈����H��{c��?�O_	|ƞx�K�R��5�K�:pX�u5�AN�s�z����`a�G�Wc�L��z�B�fM��]��̾b�8F�y��"|���������=��8�fBx������	�����r��ve�l�9ѩf^
}Va��L&O�K9=B%�}vcGCb-f�s�����G�/�HL�P��ӭ��~�l����[�z��%��zo�p��a�Λ�+�v�CS�b2��5֩�����K�դ�v��A���+x�׮����g5��`ȱc���؎(�L�Ջ��]�5�B_H�*��V=n�]	}�Lm�u�-��f�t՞��6,���a��0\��q/j�������47�?�U+C9�=��˖޻FSX��[�Ϙ���������P����О0=��[����3p"2`�b�2J���e$�Hnp}W��ݯEYȌM�l�����>�:��
X�%E�,��R���f`B���H�us�R���x_��]��Q�iA�u�F���#����ƥkS��J 
B�ύ�V��#��-�&:�-�P:W?��J<~����GmTkڮ���Z���sb�����	k8$��Ih��}8���dk �0��h,Xb'�r{u��V"Vrs9nB>���u�NGk(��^���Rº嶜�c���=��O��G9*��&5t"�Ȩ:�C���mGn?#��a�=��9����BH��R��[P�^!�p�vM�伃�D!�+���1�E2�P'PL�M�aB8�H���qB�W��E��7߳F}������IZ���ٯ<h�4�t��S�K����eulM5l� ;�Ƕ��a�C��(~���7�~)�%QF���+�{��SZf�J�>]�e�3���zU��I������.DUH�������`u΃M�ݷ�g��?���͎_8��I�BF�Gj*
V�e�%#���ʯ2�!�����o�y�oo|,s�S��1X�M�b�s�ؠ�WV	��8��K-��6c��x|Z�3�<*�m��m�l�"RJ���B#�;�颡G[���)��1��:S|��Y:��ѱߨ�b�u&�zzH2�y7����v=l�"b���-q�+r�D�ݛ\ ����md:>�r7��S.����L�5=Eͼ@�%���[��D�)��A���g��K݄H�����$Qv���lC��"�lLx�:]pk�;n>Λp��m'��U��B[�L�c��L��'�˂s�0��!�M_����/�	a���l����f�U��ޖ���sw�z�jk�͊�
�}m��7��TR���iѭ��D�-&�^��ȡ�ۜ3�,ߙY%����ƨ�g��mB�N��	�A�� ќ$!TsB-�PE%߫��tStU<Ǥ��UD�i��H*RlhL`yc��/?�0.(���oSZ�W{C���e��,<�zsSQG���
z(w�t!ݯ��+�-]�Re�:���}h�T�P���]r�����b�g1��n�i����{>�I���Ú�9�y���Q�Ԗ��f�\�k���H!�y��1n��ǝ���Cϣ���j��U��0�:,G'�l�4��뿹J��K3�\����{������Q*f��F~�fgɐ�?`W4�d��P�E�C�~>�謊�f�h	3��Q
� ��W��E�]�-n[5E@����(�I�Cg���&���=�֕�S$R�O����.��O�e��k�RW��IPm� �X������U"
��8fh�:�v^�q��3�-�ֹ�Isܣd�0�׫3��q�?�@9��Ek-�����QS0�jzͦ�=㫐j��u���jf0v�a'ʧ��g��zi��a��1���={��X��b�igE[�+(��fΆ��~AY�����:�W�	� �@���{y���95���ӷ���γ+�>8'];����f1�p�T�^��>��2\nw���}
��G��]�l�����g���Z�Qm�1���ARC�T�:���c>�P���Ƭ�T)�@�G��y��1`XX����nB[��%k��Gi�%H����]�D
�'���:m�����2�ܬ�S��6P����V�t�h�n�'�o$��y\
�b �}UҚQԉP�~ɣ�/mk���>�Α��������PD�X��(RY���d��|g�ゝ��\|�c���$	���|���C�����1�*��_���ky�����Z�cyK��/Z��H/��N�W���$��/א��V}���ay%��Z�;�Ey�ڊ��¹'+v�{��~NA���B� Wiv��̾����x	Dا���K�b�w�'�bh`��r���d��������a�A�����=���UI���,�7sS�A���"2`��؍kGmN�9�w����U1n��߬v�[�N��3�b�X��e�:���el�>��2��=��-�&��T���	��;�P���H�s�h4�N�� ق�q�ZD�{��� Z��w]n��;ӗ�l�6<,��BY���| [O�σ�����D��Ξ��OI� �4��zڬ�t���Ş�.񌂗L��T��oZ9�	�G��z͉���y)�S͆	��j��?��g�<QZ�e�9�����L�Gs��w�56ٕ��O��brK����{��?4�w�(�m]��02t���d���G�]�f�~�c�T��U�W��O:��u���ݾ�w��?���ʿ�cճ����W����2¾�B��05�	�xV�����z���NzJ��>rq�	F�Q5)�����Ѧ�lO���j9�?D��__��ڛ�K��]�]
��."��h��mP�\�Z>M�D���5�]U��-�"���F��
�G�&�W[�y��r3�a�	 #��*O�d��:O,~'ݭ�R���cV�E����e� _NQ���X�s�~�a�;�e��7�����O|q�W˿����vNщv=�I备W�8c��h��Oڭ���ft8P�U��|d[���-BpT���m��b�rY�#�����S�����6|���Dta�	�Y��@�#�0�Zc#w9�_j�Ȅ�/�ݚ�ݓ��t.�i�&ܠg�Ie��q������y�:*�h���R�W,�<���+��\8�˃�U]��̟H'8(�^�(H���j#�^�2(�� i�G��<���x�#�����7gE	�x���(Ah�K徉�v�ڥ?�m=� �L��L�S�#��q�\����RI�le�y� 9@~�6s���}V^ύ�l@ݩ�ͫf����	@򴪷�|�lJ�3=.]Iɧ�������pB�����8��v��pj������?��O���7(�Bcr��y_Q��{���k�~{	���>���U��t7�N!m?M*M/����bR�%��<��L<�=Z-NR��.rǂH�h��"9
&Y�����@?���]3V4/��c>��oZč�r ���.�(:�� ��A�kw}24�H{��7<��3V���:i��]/�Z��N?)�_WL�2�T?�j��{� }D�vR����U�^�	���a�4��y�^��	(���)1��_Z�%�����[/�;�'� �H��]��H���+4�h�����"��sɸ�$X�R�]'��3E����scU�uk�W}��m�6@`�ʷg��v9��E�k��ݛK�=�Ǭ��h]p"�D8 ��y����]��ڬ�jZ��em��������Īeϔ�B)uPCFS����d?�Vwm�fH�g[g�̌�1V�b��w�~S4&�L�@b�[�V'�i�(��y�9��Bd!��x���a��l&*aq��ڹ,�CqQU�z��%BK7O��r~���/L�M�%O�<�a� ^�����6��F}�p۳i���O�x��Ɋ��eF���S����1���	_B�
�*Y E��n�����C]����e�����{z�ʪ��j���5^�G��+����㲱�מ�~ќ�0�˨�ql�'JsUq���O�k@"f�$d&��4��I@�K�H??�`��W�y8�� �����ER|$}&:���[�e�CDHغ��j�E��f�y2:p����5'��܊HeQA���ӧD��)���Bʷl)~v��*���.l?��&�`w{��0=��O��~d|����,j�\�e˘�6n,�﷤ٙ���t��ҳ���wT^y\ޙ��G{���Ҩ^�Z;�P��z���8%��M$��T���%�U]BL�d9�;����_�iIR�'n���`���F��'�t��� p����#�St�.�՗��:$46S���I7�?08�A~	uBA�)8��<�M�B2�D�" ������go��@�!���U��.`��93"�e�=Y�(�䪍�&|$����ŋ'̞\`Eъ���Ί���t>e��+U\b!��Yxw3��P��d����I\<���m�l�~�Ԫ�`��*�3���-2���Ec����*掝я����;?~�7�����o�ض��:C����@�z�dw�S��:+�\���T����6v�UT+x\������Pcq�ɮԂI�\�[L$�AM�P�.ۉ�X��Vi|O+^��/�a���i4�B ���k�{H����.��`���H�^��������\&Bq;�.�xoJ\9��w�t<A��/�Y�~�䖅�Bi���X��VU��V材
V�xg����Dm��"��)�����S� �3�L���H�l�-� ރ�X��6r5(�5�F��yR��N�F*MΫ���o��UA{?���sD���$KȆ��f05#���3\b	�E�
"*�\�<��XdX+��:Ṕ�9�J�2o�b�;��G�R/s���
~1�p#{�U�kȀ��A��~Ø1Qr�I&ŧ$_��1��3"�]>���J�
W��$k0A�Z�I5��G:���]C� B��Wl[��2�a~`�Sy��&gK����	@ɦ��.����~@h-�D�*ᝓ��: CE�j�{��J���V-6e��@U�%�e�#�C�y-�Z�����+ϓ�������/Z��n��t։=3H.3�&2�/�5P��`��c{'�*�t.*h&j�G*�Y{�N�R�$�^W(��C��B`�9�񒸤iI���qcG
��U:qK�_"zh��DT�TyG&���m/f�Y��q�oY��&{	/����.Vbn�'��ת�;)�o��FgX��Е�	�s�?�Cg©'�(���G�Wj(rAQ���;o�U�lt�����&��E^ԛM`S0�'!����c��Ǡ��*o�L�.} CN�����tU�S�0#o�4����lٮ/OcAܩ�6�w#`s�������N8���{Oש�P���e�gN��|Cvބj�l':�I(�UK���s�9��`��t�֍pF܌ī#$l�_ށ�Ņ��H�ul*�>��/i-�|�py��s���<����
̸�Q.�-�\�㍮����~u��c]XY���
��AMM�eu��᥷���+����ޓ@����'K�.�@������魐�$ƽ;�y�ju�R/�	?��G�g�g�N��h�G��7��.:D�%�TelC)Cz�����NF#|�ˎ�#���1��C/-�����u1�M'��xN.�v�� �C
�'�>M�YW"*,$��y)�:x�ٮ��/l��
MO#����6Ϥ��#\n�<��b�+�¶i:X��� ʷ�4rT^�	�3Sܖ�Q.��^Hު���W�j����С�~�	p���]��5�C��"ߜA�M���;օ�x�&]S��H��a����b��'�Cb4�*��%�R���AV="�ɚ�!6�Kaf=׬���z�*@]�w[Θ��DW���T�7���76#�١QE�����E�]�z�4�Ͼ�X K�B���R[��g�jV��S����+t<�[�L���ᩭ���/��bX���HD�"���-��f����,����� ����'�:��v��Րm�ܞ#�K��a�j1�~�h����"� -�?|p��v���d���IWͶ��ǅ��ʫLo��!����P۟����ё���:�����J����j�gm�"�V{��7��{mzLX)q͵ml&2�˺�ٔ/�4��5)��b+o'�cB�G���
^u�m ��&,��3^Z}����t��j�8|Q�a��/j�.��&�ͦE/��T�y�!#"���7���{���/�܎ھ{/VpmQVI�;.����L�_�J���<w���,vG��)<Jdp�������n;����؆ ��[fݥ�X�U���> ��\���m��􌭕����J�����!��<ִ�}�qݻ��C�,���x���x0�V]�J4����|�Σ�4{#O�(@�G����-��'�/=Ժ
�"v��¤O�c���a��[��@W��s��!�eKim.zyx�?�q"��?�CV��C�0gd�1�[�����	�:C~�Z�%'�2�АT����J"��sH�r6e�;lS_:�e�5�p� �tY9�To����3��{r���]�/��W�9���K�&#R�Pގ4>+�@K�n�=�)N��r����&����.�Qet�n��ςcI������M��֠������o�Jk�K[[���b34<%�^��a�5��r!��(g5�BS��P������`aA���~�!�8�ó�wײN֮�;���V��n�lba�3�ֻ���A�������9u.8����t�`���&Φ�zp{w0S+��,ļ��p�K�FlIUy�i��0ۙ��o�sWk�kZ1	��PM�Q��˷Xn��x�W���4�x,���6{"��'k�S{L��C-��&IK������QZ�@[�g����s�KKPD.`w&`���)Q�8�=�6��㪾�NQ�|��w��N����>���vpـx��
� nF�Ө��~������@.죟	�x�w/c�&�1�-��!|h��_���v��������񣳑6���������r)`d�T�G�����bH��	J��pL�Z�\o!zWq�o��~F�ď1"0"+�:)�Hv���6k:L�ޟ]q������W*Sw�-,/L^[(MeF2�`x��BkY$;$�����~��{!��up�࢑���:
�R;H��J݁��W7�pt���ھ�����y�:Q9�>���9���� 0���O8$p�v����@�O��'N<ں�^�,N̡X����=���I�rMs����M��9�1X�zm[��CJN��w�,�6�>?���HK�q�آ����Y��h�K_	md�7ʤZ.��]����"SSx��Ţ��W��m
jϕ(���=���V��<���s����.D$��vڌ�NQ!-�d�ʭ׌R��m^gd�L��3� n;�㳇�N
�U8�H� �F+���<[Y�G���3A�y��~�}EW���b[�ݳ��5�,��絭2G\�<3�]�����t帲�+��ba&�:o
*/V6D�['�u�j�����˿8M��{���녤��f~O��m��=1����J/F���֨ޗ`V�����Q�/MǮ�dͥ�I��4!�3���y3��:��!c��RZ��]a��`��bBeb�!�q�+�n��o��:B
Y��H5l��\"/��a{j�J'��
ϰXJ��^c-Ф�_A�'{�{�D�p������.����bf��4F%f���ϲ����r=�7���r�D����=��1P��=�P$���B-�s)K�]�f�T�O��y��4]\U2�Eڵ@����D���5�S?]᮴�f�ɘtCEi��
��q��:�a��4ڙ#ӧ/���Lt����/n6�;`ݔ5�9�B��kz:�_� I����N*�<,{댖�X�2� ����t�J{9p��٘���v�e�<���\f¬hR��#3���`3^�����K}��+Pj���"h�L�OYDꝅ�J�'#@��T�%K�~��]�?�C��w!:�3��q��0��~�UF[B��z�8k5�f@r�A�r�/�FU9��Ѭ��F��50n�g�S٥�=��N��y~�P�V�k���m?D�l%���ʦ��i�VpI�x��0�Mt����WM��� {��aC��|�t,X���p���M�ހ�W��X!�U�K1�����',f�]�}�x��YK޹���6�Z��Ʈ�������|��a��K6?=���Y[�i��� ��E.�_c_B�Fx���\��c�:�H�!���HÏJw���2T�&�z��O~
�=��"��G�ϙ'�&������|�gJ΅��muwצ~�+���b�̚%`_3S<���1'I-f�tJ^&�ef�E���U+��� �R� ��5�s��Dzɬ�7��dF^Q	ɜ��&դ%�������P�s�slo�!/*�}�J8P~̦'�z�<oRd�*�<X�l�V��%�ycz��X�OTuv ���Q&�����}��q���4<r��� H�.	�$�n ���g�W��mnm���	�j=1�����L\�1[J��udL��W�R�3��Ƙ��V���Y��|����hOV�fR4�9��M�	5"Q �CT�5�t��r\3�b��ל�l��� ,�L�[��M�c)\�q�UԆ�wv��)= \�0��enW������k1�	GT�<�@7���;�;:j���)���\�&K�M��	� Ռ'C\�2��ߗ����q�N���g�S�[�n��H��uAnbs2_+��@�S��o��++��d��·�Q^�Ҝ���mH��fsF�I�22~�ϱ�C�t���:z���ZyQa��7�!/��9����`$�$S�kv�W�&��f�K
�J��U�9i�>i�g���t�I[�����F���a^J��W7'u�r�	
����c��*7Op\n&۪~��
;�*�K�v�5,�8���2�� õ��Qн�z��,���L�]\Ud��>n�;�L�o�Tdm��r��=��aL�����ne<8�_��!�T)A��ԯ�v���5�����	`�bK��!�Dg�������)��P?�r�R���1,p=���O�3�f���}���� J(�������Nd�C�[A⚁�@b�'IA���8SPM������5������ϩ��Ā�%�WD�C������F��L��q���0۟$�2k��é�7��_;~f��*�#h���-����P��_�š��l�FI�~=�dԯ�%�p˿������2����*�x��I������F|��~����gYT{>�CQ|���ܟ�_��d���%bQ��������aY%آϮ��Fk��'����HX�5�������[���U�-퓈��^�>I�Z�bJ��4��0l�q�WW����v��O�+�w�WV�pz�Z��w(o?�x�p��m���}oFnSΒ��z�I�L�6D��b�9������j v�k���A��,Y��V]�|�}qꊬ͡1Kk
�?�_���R}A����لP(%��fT�i��-d&Bc�gX�i��w_�.Y|��tq;�S�8�UiQ�=�,�[Rb�A�'d�)ZN�(�, h�Y�$��#��slt���5m�����#;����>�,�H�;��k�R ����T��E��)����:gaزzcf�ο��An
��Y��	��`�ə$�7���}�iO��Me��Ѐ��~����).z����WDW@��]~��׫��:6Dx�@�*��+a��"�U<�<G��}3�&�x��Λr�c�kQnsV��KI����}�c��.r�v�s�QބKXut��"�s� B�aX�T�d�}��s�����=`�poF\Em���L >�����4+��iQd���O&�'N&:���g�Ҁ;yܢG�R��<`��j�F)���Ec�MP��.���~T\L�_.ˢ�=������vd�=	��WVKx�����0��=SB�o�N�]��!5��.��Ȇs[�����Ħ�H��7�k�{M,�'��@��.s�c��rQZ���%�ZnG#����a�_U?��2�H�"�N��b����&���xGP@
i���U̬�'��?(��kD	�vq_FVPU�������V9P�H�%1-��\�[���,�!�b���~��N�%��݃�"]\%�kd���^:4цm�_U���"'��]�E@hu`b��}�yzB��O�c���Ҥmd|�~�"��j��E�����}Im�B�Loz�O�U��g�>�̈wx�����O�J!ZĦ�~Z=�"%Y�x�?v1����d�<n��Ekx���҄��{F9L>V׽�Mh 0r@ߍ�$|�ȍJhR��������c�[�hS��»~h�0�6������mPUȰR_�N�'��k�8)�be����΍@�A\၁���뷁�a ���U���
Z�#3{V��C=j�E.~է�*L��%V�+�̗(Qͭ,5�
��o��Z������9]"MX�2�;�9�F64�d��'s����V��اht� F�>���m��0�&d�ހݤVCˬ)Z�Z�;V"���[�כ�)��߸���97|�xN��8�׳�/Q�#�밂�}�¡^�TW;9{����R�C��P��J8F�9��3e�q�/�=&�k�f�&#�����R�wn��ݖ������.?�q@gH�X�d��L\��o<{��,�SA�Wm=W����0�BZ7a�����'�N�s�������,�b���W����J��5a��1���H'���˨�t	aWH��r^V�Fz�?�)a�����y]@���<d�/����d(C!�*Ym['�-���S�Bd�,D���.��D?��6�PF����[�A�ę9��´EA�U��1lF�Ô�}Qx��!J��z<�Z�2Q4���n[�'���yB�m�}G pkn��N��g�C"�)׳z�y8~���'Kw+�u�=]
��u�xh~�ٵ0��tCw_�.G��}u���k$���}�l�_C�<(�^�[�<b��j�
�P[	�'�"w���1�8�IO����*/���� �)�f�h�t,�)�ӣ'cM.&�ϕ��.�",8�!��L>�P�d���8=�l�EO���'y`t��6޻��b�9;�Y~	ˎ�<��2��|�I��Փ�]��5�j=/��#�ܘ�K}ݩlOsR@ʩ��z�l�	��%+��@�e49u�t��Q�ًW��P�p�;��vƌc: ㇍�a��Xk-�ѻس*
�e�ō�����B�dkb���à�c��k��E{�A�����m��W�v�QP���X0��)[=_7i7�]N��Ӥ}��`�iE���1\��wO����a����ޚ�Ю���
�$�rf�WJ
�qx��>�El@�*\!�N�W�� �R�
�H��4�]O;ގ�D ��=��}y�v
�@߬E�LB��&Dd1���s-��D�l�kp�uQN�����Ű��tH�Iq�]=%x;>�V�b�v8[v���o�4`+0d2w>c�j�|ޟ�Bת�H�*0�!�������� ަdM�Ξ_�*2��o'w�)�D8@"�<@F;�զ@P��"̹�^J��G�T�Ʉ�78���3������.I�g���yQ5�]_g�Λp$�;j��	f	��ީ[��>>T��з�1Dt#l�1[�0B�Z�B��8j@k���F�G��,��[�B��Y-g�b����<)d �fU?kߕ�>�v|U%I�����ˬ�
h�V���*'�L�M8�g��6J>f�jܱ��	�x��`uciMm�^8�-��,��#4�fB�8eÁ������E*\\Z|ځ�{X7��a������"Bl�c�F����T����c�}�q|��j6܁
�o��Ģ��+�-�Qfꉰg��5.ch�{���]��P]�Qq�����{��EB�,�.:,G~�D��"XJ�_�> 5�z8��T�j�/�QD'����*UE%�ƕ�^ai�4Mj8�]Q����z)�ux��\-��+�=��x�x�����Oĩ'�k+6����w&�Oi���h���fQ���hl8��kO\�����3S�t�'2[$��v�1�ĳ|�R��`�����sϒ��O�L��^@!���7w�n�<C�9��?�\���Ul[��A�uwMD;E�wԭLrH�!����x)Rc��D6�_Rε�r�]^p#�N/[�%<6V��R�t\삕]��#˃&�-�*�i׏����֪��D��� 5����҂Ĕ�Y�>1�a�:��E�Yo-��Y���!I��N (5��'E��$iAV��Ց83�_:>s�Ĥk5@tR�l�[�����(s����/|��� �:]�t]�^p
�줥ˮX��L���j�R��p��ßc���3n2 �D~�H��ٻ��1D?�ƻE��0��u���oA��(�)����"�+�Z�wС?:ţAy誕���ߎ�g 53l7Z��3n"B��Ӆr��EyK�,�H����}��Y)���+��G(��i�-ܫ�8'�	��0߉���``uE��O�0��$��gK��7xG�� *��b�7��UU��s@4�>�e�>D�Doo��/8����τE���!;Pm$G�a��y&\<*$m��^c?;"rk�,��4(�dpi[<eaf��G���4c6��6;>2��^U��u�4��Or[���u�0�-�Al2��˛��H8�F֬EdF�)�ܹ?O�������g��|HOY�?��+��j���S��r�\�\�-"]�~ ����o�4v�b�M0���Y�����N��tv"Z��c�����'��;V�˃k+֢�v��1��`[`�)\,�xv"�'4l��;����7Ժ�g� v>e��!x3�c��t�����+)�͜��<�E���>&�;�Rf����#]ǣ��wS��n�q:"�}@AW�V����-�xB7��Z�A)��Ï�Z��P�*�>�N�J�)9A��2U����%Ǌ�Ń�[E��9�W��E�!�V�0lR_}����	���6�bgf��9ebQ?H1����U!��css��H���3b�`Q{dL[���bx�|*�~2����`����m����@��X[�������^A���Mg��֋)�ȓ�1i�&�!	��]A�U���B|�,��^3�-�5��И���fiG_���7����p����]��>��/h>����1x|8��\e�����T�JGX�V��0����Z�V��S5����E��7��| f��S��%Vz�2*3�7S�\O�\�#e����Q�c�����N�-�}k�u&���N3��g4�%��,�����p�DeXd�1�n���${��M9�q2���1+c���^�p���`����@^N��i��[�HvtKq�2d�LюS��뎩�� �$)��fϿ��G �.��^~�3*g�;���C���(�L3�s�M��Hz@�!a��[�@"�lm:��L�l^&x~̭�M?e�@��T/M"��~��A������+@�ԩq�����/�O�RѠd8Yx���(q��i\ƭ�1�'��կ��c�3Ɏ�)Qs���!HL�q��ϗ��j��g�c	%�K���
6��QED��5��r���������E�;�3f�_�1�!����v�@�U��4���w�DhCf#��}��x7�P^���.�z��{[VP���E�^�m]��6�&�tYs=[����A`��z�.@��3m��1g-!hy����b��siJ'�BG�<��;�E�������r�3 ��Η1�����4��xZ�}D��;L��Р��!Ţ�`O�����jl�����ۤ8�9krһ�:�[ ��q`�O�Y]�9�Ѹ@~D
��եb(�� �@��߳#
�~F���/�^��U(�4���!�]�-5>���� �T��m���Wh�����

���0v�>M2�t��$��\�
��ęW.#���sL�՜@�_xz����B����w&���1��A���ш���eE7��,W�����q�]E��7��<t37{1��.8�Q�E3��h.��:\r�<�~�
,b=�X̀׋�j�Xf�ws�W�$ˈ�TD���3�CN��R�mJdfb�f2s'�C�Y~�)���'�{;��b���s���M��B:�e&���&g#�:�q΍�G|!���Vb��	i�����rQ���)e�ܾt�'d��ɸ�T��\yY���:g�(lŠ�pJOz��p��Hi!ٲ�'uj��`:�B��/����س�cM:��ܹ�O�1���'��)�����������D����!5V:�m�פ;���L9��18["��� �Ͻ�n�Q��ۭc�������hյ���uOR3S��B���~��|���0! �L(�_K���Z���c$b�o9Û/Lv�E0ΕMѣgi��wXĊ>j�6,�e�nUs��a���j�� MA� �+��BF�j�s�`�^�;���8�1!s��	�ײ��{�L7d��L��ͬ��X���
���:�(�L��Bn��}}Id�a4����Y���_��+�i|��.���|nL�������?�Ak#�B��ܲf?�A��O	7Iſ�M
�H�.5 �yW�3��a�{e��������`�qGn��=Ͼk{��G+���	>�����z���w\�?��0DG����x&����"Z�ݍ�����Qj��O��RW����s/!�W�3���+��0/�Y���W������{_ݔ����5̌~^z}`] �W:΀�+/��!�c��@ʮ`[��R�c��+1�������D� �C��k��^w�nu^��XXfeп���*�xO�ջ�a+�z���׊�b̉��"��X)��^��l�i���.��#�j�<N5C��G�>�p����3e��d��n#(����.~�HX��ͦ�=Yg���}��	Y�������4~��Bt�R$��/T\U�4h�@�����T�0����I\a\E�W�����I�HY��00�>�s�nu+��B�r8����+gI֘ӏ1�=c!���A����q��u�a���M�n�u.��1��>8jvi��`ߛ�X�F�uo\��wu]���(�k�c&��Ǣ̻.d�����kx��/r��Z�M� �!�a�H�Aǹ����/�<�mf�k�\+ѵ�o��Z� �l�����ؕGhW����Ӑc���˖���wha4�))�?��D�c�=�7I^ ����$�R���:E;Q��O"</ؼXs$�R�����/��ˎ���g�`p�"ݳJ��g��Z1�(�L�\g_bC��<�o���K�&Q9�Jb�a�)�0�� 1a�gF]�Oyw��&�z���R���)���U@������oz�&XM�������SmioI��v:H+����ypۂ2&��t�^pM�{�=���K(Zi�)\�'>��
I `�1n�D����:'�g���'r�I��	q z)�{��m*���6�-�����q?`i�c���J�/��#�:���&��PDo+�q$� �����t?���z�P����̐7�҇�meK�����y�P�$���9��-�O�]�}�Xm{X�kEh<q�q[��PZx��#�0�����X�	
+�x�*��P�Z|�����kY��F1X���P{eu6�(14���Y���@c�/6|s5�v�)�����O$�^r�tyz�1��d�J���c�����J-ǦV��Ƀ��v-O�����,$m�h�����W>�(0���̐~-����D���>L����Be�ҢH��%:�F/��r@�+�oW���orHĀ��2T�χ�wY��ї�Y�c�$y&L���y�����&r
�V�m �+�����V�	6ß��m��K<�x�Y\�J]�7�Ƅ�q��e��Mr9����j��_�/N��q���\�#��ͦg�^H�%�ڂ(G�|����O�Cbp)pW
`�.:HN�N������Cl��%�*,�\~�z�1-#��v^sL{SF��ZI���f�u���V7 cA����օZEp`KuS��
^���)��T0����A�4�)U;��F=s���Bw-u�2'
�;��ߜ�ô7��_���hJE�6�w�pJ���u/���~��\y�>�9���x*wq�� _u�C�p�\<�tvm���N�C�d-���B^<���u�#�A��L�o��Gƚ�ҨԖ�vipR�+/����Pi!zi��s��Bݒ\�٠`��s�M�D~8�����������\����V�U�KS�շ��'�:��6p�,\r��W���.�2��uۋab�e�#XZ��yxY��1T8���D����Y��o�����D`$��� ��$�0?z=�W���Z����cL7��4���dn�1Zv�2���0x�-�D����84֦C���͹�=X��� V-�-u���|��˒�V�6���JR#B��c�V��#��v�4�9�����p��i6T��\u`�n�up^m<%?�Oe� .w���[B�d{�QE�^i5&�2Y� >�`��-�+kÃ�������Je
��~1�u�x��עw�|���*�l4�>P�"0�҅�6��)|c�[b�.{�&��k�����}��eZ�q�׵�X������Q�Ǌ00v,����ݨ��k/Hcb��q�w����h@�g?�\��Q�@#�i��]$i��{�'�
K�e�y}H�yZɼ�;��%�hc�-��I5F+��(�@���cE*G�E�L:��U�.��`�k^�O�%k���OFZ !`�ZַNa䤫���B��}ܣQ���)��8K�)�P Q�hz��'�0W���#�]���X����K�^;�4�	�{i$6�����"C ��԰X�w��-"Y1ÅMi^�CĬ׹��v]v�ge�1ng�1��l�E���ъڢ���td,�Hݗ�jM���BGV� ��;N�}��F�Ӎ���:��n��峽�ڱ�DQ�C]��|���&8 �<��@��k���~<h�X�f_dY���� �����F�}��)Uk=j�B�@-�:oi�U�Hp���5�������j��ê �YGP�(X��Jd�0�Y�l��G�D9�L���������m��zʎ�gy z��$sx�D��ܯy�
f�`V�m���K2ex`{���0��fSZT��� ��c��͝m{������+�G]y�ɥ�1���uPX/6y5�EڅD4� r�Q�G�Lڷ���ݒV��C��PM�Ζ[�~Va�(
��+>��ac7k�ه
���^�)G�G�9ɬ�3v7g�7Bc�H��m�*OL�W��f�Uu�?�!�D�)��QsF"Si�q����̈́���G��s������hF{�_�/� ~^E�s���[��:w9�[��!�������]*�)�Nz����r��<O?�=�~����K�U��6����^'��a�t�پ��͖n��0�^
�}��֝�O�=HK9�
��B���ޮ��]H ����[�p���.jgi
E�s�(�Z���Q%���4۴�8�Wb�D¤u��^�3�[�6E}����{��4�<+� +�1?U:��ڳj|p^G3Ƀ��q�(��Ek:.���T����x��gB��4�:�V�h��n��%�4i�.�@+xṅ�T���:Ȭ��)���c,/bZ*j��yW8��G\Sh�U�L���<>5�d$'�}h���چ� :ξ��h�磉T�a��LPM��Dk�Ŧp�:�U��NE\SG�~���~rB�K��F:��^����R(ʐ�ƨ$o�6����zٲ+i#�u�������H.�H|����ĚR��lJq�Mᷩ|+�$ ʹ<�:s��]����e�������z���Fv�I諫��D�8�_:�/�ċ�Kݜ�f:!�^|���~r2 �ɐ�Z�7�W�C�y֜J���_'�6�^�㓼��d��8�;>��+��m��t��'@���ȦwG�^���;?N�����G�0���`[O��ZF����R��[.��.�,M�Y���L�����A�B ������1<g=
ʎ���,��H�eG��Ai�~�,�W���[��!��hf,'�/oa�b�j�#��v���'�$aۘ��^<O��K�)�}��x����ft�^T��ۿ����P��Nvo~۞.�R6�v��dM�QM��놦�=F� Π���>? Z�<�|?��'�IA�H-����h�I����[�*M �"mFf ��#���&Z��2��U�_����O�7�"�����P=���G�Ӑ�\��á��qd����sDK����_~c���_ �fqW�#���N��"xIk�+3�nI��e�m��v���Eup��ҽ�꿾��`%��[�Ņ�Hm���,�9���Y��©��$� y��&ca\�^�_�><�b_�#zA��b�0h`@�G�cȱ!|"��x���UFU,3�|q�����د�F��Z�5��]bǀU�}�����Ud�U|�0���n�(�z���]2��kf�CF-�:(�(R�ӯ�j�1����L�7�_u8?s�[�����5i�Ĕ����aT1�P����z��;����c��3||K	�ݙ�Y����g<���6M�Tu�Kf��!�E))zj6�yQ��Uut��j'���7��
��7���sR��.��&��ܰK�d}T ���P�
\5�7��O'��&צ�۵ޭ��Yw��8:U���RWw�ŕ��W��3��v�vԇAAx�M˄�� cfK�D�4'H�/+_W1X:�Ƕ����R�<�$�]=!+{��4�.A�,���PM�к8�쬞�j[`�#ȶ�c�^�yp��ݰ�����,�H�AJ�h��?M�pV�I	4��4\z���K�!I`FՈ�����T�w�I��Gj�����X8��bm�.����A�Gϴ�������Ȃ�A��i�F6�Z�ƨL��w������켞1?b_�A��
��;��l�2��Qa�;����r�Hg��i$���� ��"z�u7l�������H��Ck������%��<�r�Dʽ�/�X��3���7�Es�귏�x.�9I�h��0* ����.wV��.�{���T����}�pN��'�z/P+�$���&��q�4�ס�x4К>������3�.Ï����E%$��5��K3}���'ERtR������n�3�z)y��</�j!:���Ȯ�$�N<���qsb���x����H��@��6��s��ܩܓW����\�<�7�ҼA8~PiaY�&�0�}�M^]�z�L���Q�f�lN��^�7����I߿��Z��~����~x�Fyq��i-ф��m� �""?���-$�*��(�`��lx��FQ��ˍ��M)w��o��9����$��0��/�$�7\��y�?�����'�,u�U�6��0ӷ��W�{^�+H�����V0�_Y�]���N�/��W�-@P�,�>@�Q��р1Cm"x:2�8F*��W�PpTxH�[�@��7<�zw�B'�-=�����[L��]���X���zs�;�l��UmGG�X_:��D�o��B�(�z�L����Ȏˇ"���#�^b�
���$��M���̤���^�l*�M%3h �°@R��T�G7_t������D���K"2u��f��Ѷ��b�<��+@��R�� b'��P�졀�h��&It6O��i��}�1m��J��3���#�iL�KȨ��h}�Ҙ���%-PK�*�OG}U�	�l�t�KΑȽ=��"_3���г�h��Է1�NI#�a[Y���]4�TMă�Шg� e0�*��aЄK ���_BB~l2_���I6=�|6&e~Z�r���׃{�}�.�Q�d��a��K�fPMO{e5�R��E�E�M��&I[��#r���U���^H�_�w![�d�:�~�*/��M�Ӂ\�2�, �t�:�L�����fL�rW�h����>e,��/���`�1a�/�ף�#����~g���}5�M�K:�T�U��c�oy@P.N�6Y�Ry�'Da�/�.�Ĳ���y�Rj�]c�6�}�&Ÿ�<���%톀�������w��0eQ�Lx�Z��q��� $dq���q��r�{�X]5�P��~� |Y=������[�D^;(���6�d�K�������^")�7��\�7W�K���/���˕<yIX�^�n�w��U��4�" ��N�tW�e�<�h������ʟ�����H��O����=T�4�Ҍ�Y�<ڑ/m�ʖ^ѥ3e#y)�f]Y;v_b�R:�D�����YN�ou��+>J���Q0HZ���%va�쎩����,����( �3��UG�Z���!+���O`��س�ZF�#�A�l��o^��.��xr��o�-ƍt!�=!�S�۱g� �X6�yml��w|v����N��1�����F�vʐפ�6
 ��Y$N��b��d����$�~��@V�8G������gk�L��jk5R֠M��-��N���gF&gx�z�n��D��e�� P1U���A���;4��8���Z}`E� �M1V��f�~�!cs�~��0����o�;��;-%ihdNUP����Y�?�T8b�:Iډ{a�O�͏�r`dAG����N���1�٣L��;����ӫ�ZP}bD<t\�_̢aP�����pXX�־-�V��;�
�*���Nv�Ix?��]��Fy����'R�D��	hР�欥r�6���s��k��(���o��.#�}���/+��h���pp-uB�.����}~x J��MIN���(��	f��͘�F���t������I���:�"���L�h(��L`�&�<��#�m�$���{S,�B|�ݬ>HyeDՑ-G�(��4‰�j�D����Z;��ݮ�2&RH6��ޞ慓�Y31�!1�àg���5��A~��b�j�\�0֔�rǨq�ϿI�ő��c\|��Zfڲ��>�}iz�4' ���h�	F ���.'��
Q�U�7vd��&��(�G�@�"E�X.Tq�tC��KZO#m�/ʿ���-*)UuJ���n;�8y���Em,M7��sqnȫpG�Q�hy-�A!���/EZ���H��M% ڼ�۵�K��׿�ǀ
�&���-}�b��oR�-���a�UFr���l��l�b�aClC0pu�<g"l��k�eH�N� �٬��1��j�pՆ"�5�W�&�V׸��#$Wv�	n��k�OYm��V�5�o
^-�X$.)!�ZM�Mg{��0����.�񕄶���Ϥ�HV���c{�)��'6t���?�p�S�������@}��:;bNZ&p�# ��|���(8����u61�� A~����f�;J����郄���%/_�j0�̔j�&�oc�Ϊ ^>jDDS�j�R�^���)R���J|/%:Ϫ������<�[�o��e�*���W�e_���2�3��띵w���-���_�T�9W�h�e��[K {����zZO���K03�Š�W����_��X8�@���Ln�{3�Q�$"�0�\��l)���VMɦ�>��Ar	Am'NJp`�_��+�E�ma�\���\�Vy�v�>elX����B���N]d�Xݖ!GM���6[*0�ʨE���j݆	�/�-ɶg�O������	�HP��m�;k��s 3�-��f�D7��)�{'�t��z��]p��*���J��*���U6$�~\��`���u�=����,~d��9��q3��� 'i�p�¤|�M���;fA8��7�5�R��F1&��˩�%K�Ҕz �FJ��uu���ow��#]Դh��d@����x��Y3<C�ϡ~7�;4�R`ͣ-1���
Q�	]Oz�r��&��.��N_����U8��������v,3vw�Y�+�3��Ƭ�[ይ�G��<�>>���G��9���8ᶗ	̐���RWY�"��|��Fy��u�����#�zPqQ��_ ��|-�3�
7W���h��[\Qkn�3'��{��y�vH�JHn4`���!}����S�ĳ��a+.���N�T��UX���g	���!���o���M8i����ֺ��������2�dWRw�\�2u�\�B�Zje��,�[)�66�����{�|���)�5�����׈ރ�D0�1��u��(a�;D�}��3�N�FyY9�fK�m-_����od�۲~F	����i��W���Ȕ���_�4��y��@�CEC��t#��Q��c��
A�m@(}��:�u �#g%��U\�	�L���*M�"F(���rytb�먶=t�:��>�'bE�@��Ѱ���o�g�\^��
��1��}ū���d6hd:wDD`�F��ԁY̖�g�P�)`����w+�Ui~&�i�@��Ǚ}�O���v��a:��5jװ`{B���v��k{�]=��-2G������p�-$�Β�n�Y��� ��
̿���q���XY����k�L�2i;����1�%�1i�w��������W��-�=�B��*)��w�L��Z�ҧ���܃.'�hd
��d�Q�`��B��G'�"���������z*�8wU�2΢^�S��D���j��$5����'��I:H�S�&y[ߚH�e������6����^�Ϥ���a~�s����Ͳ��c�=ѨqpHX�x7���[H&��C&�6��gK-3�-����\�q@}JZ���>�b�#E!XZ�SjQ�q,;?���1N�&v,��G��C�a��8�գ7�������V�1��Y�,>MM���{͓MǁW��O[=D���);As�Tre�z�c�j�mr=��x�c��T��I�&y<���O�F��4s6�eZئ�|��Ы:3�a񕡸��N�l9q�=�[#�[3���p|��bڮT�"�n6	���g��1Q>N`�p)�iY�d1�$ZCB^č��+�#�f�p�(�m � Pt���$ �%x ���㮛��pDT���k�,R���".�A���n(�sٜon�P�R�����vq��5�J�)�������Y�Ү��0� ��?�:�?�j�0ǁP�ʰx�=_��xV�sVV=&��d�DǤ׸K�����V����'y����}��(cޙ�(�����f쁷����Zj[RF
6}Hx����Ɓ��F���lt��'V+3o��-�eŠ@b#��4HB�<�^�l�����E��=��q(0��#�������fk����nX�Z�2:R�J�.P��\vɖK�5�É�("���+xq�aNCg�c�b.��� ˫ߵi������-������䨘NQ�
I;�dk?$���j��ׅ"�_�Vd8/�M�;l&����4��Τ�E�_�7�X6��_{8�}zE���"DP�����k��@�h�a ���_ZV��쾚v<����˾x{�d�b�B e�L�j�7y����9����f�:O}]�򫞧\)=E��5f+1[f���܄��y'���z9T�5��L ü��9_�0����I�X��J6cW�WM������4�gA	h`�8�������a8���O�uF1�U��~,��i�["�[9F��������	��cN�7���3g�]s}�N㑖Iu�J�@	R��Lʯ&TC,��R1����S��� �UCKg����);*mZ��K�FF��6���K̓��E�5�X�s<z43<��5�͸�?��Z9ε[s�V 1U.T>\j�$_#�������;�V�6&H:8�^8a�e��k�L3"쳓�$��7h1R�y���o�{�N���I�DF��Pfᾯgg���ς���xQ��2WYl)���8�'5�����.�d/Q�"�mg���� M����7=�-�M����ޤ�PPU������em���ՍR�t��rҩ�9P�X;��v'%�d	�|x��&�Έ�P��}�LZ)�#�=ޱ�"���Oz!1��53�3���Z�d#�XL��o�'��g_��^��i�6�J_t*^�����9��G>�gTx�!�}�&kW*����R[\$��`ZTeݝ��>K��DqTP*d�۲/GJ;�Bq{��L���O;�9�Ԋ2�>�ݚ����ל�����F�l����k���3���UE��� �K��\�Nф�İsmF�[#P7P�G���m��U?�)�	� Q����V;�˿l��ZX�ML��O[L��u�W�Fl��5{�Ɲ�tm��ؼ���a��y]|;B\[8X* n@N�B�yv:*xʐL�R����ۇjb���Rv���6��4+.�-�j~���>��V�K(Lnb��x”��Rn5`�W�D��Gڲ64��7Q�c|	��hmpp�fioOc-�O�U�����z�tﵟ���{MD�G5��l�y,&�)���E��{Tt���О9�~/I=��2��mN�@(�l�%�?өTU@��IEZa�l�¤�>�ZI��F���Sǝ��^�	��A��sHj>���J
*�� ѰV�17�7�$����#2<�J�-��V�m*k��`��E��U*v�Y�ׄO#�J?3I���v8�CE���:9r;K��F�W�����j��6�`EZ���|bˈ~ʧ�l������Χ�D6g��"��I�Wa�?����D5Tj}��Ɗd�}/�[b�ٕA͞]��.�����1Ԛ�#�S�p/�ϑ�!�6Zw�*�ck�Ȼ�t`� .~<���;�"��o��#A�؋������Qtp���[��Lw�� ��/9��+<b@��������2�&�Rk�`�E�E�oi`�g)�ND�;:�^S߮��?u��U�3br�y�E��c��p��H��$�u��W�b|HC�<�笜j�2����K�p����#h�X���C�|j?�k@�2HZ2%��iS.��`$�K��_V�٭N�k%_��\b_��Y	:[�$pw���oa��W�Kt�O	���.U��&���A^�X�������*�B��#���&E�mۡ�9�7q�F�W����>&�U/.�E��t�x��h0���}P���՗��bs���O��ЮB�s�-�v�
��,��`�ԥ��:Ҍ�U���zĸ�׃�-�s�+/�\(3]��=5�hK*|�Ov��p��F><���=�n@>�7^��M0䮄��F�4���KL@ ���Mx���0r_=v0�N|׹x�PO�;��9 t\��%k�<B5SiĢ�>fi4&l��)��a$�Ǿ��9�f�6�X�G�╋k��K�W��
�LB�����H|����EP�{
�R��w8�؍Z���&�z3Ó�Q>�p���M��ROP8�)�_az��l:yW��LI �EhI<�oZL����HQ�	;:��Fz�zf��xN�G�V�ł�
���eib�#n�������黓�2����sb����g��[>�����_�d<Ĕ�I����c��q�j[����\?�B�Ȭ����3E��z�[�W��Љx��|�>|b>��  7�������ᄲ(9�\ٹ�6~0��Bٛg�v4�P�L��НRn��	^�q�h�S��ItXǊ��t&�;?������`�L"`Ⱦ̠��q��.'��ǀ�L5�4�5�n��1��<�����k�Uh��6q����$�E̖M�������6z�?+���'��7E�?0��*�
�Y��C�$i*�G�*N'6�g�i�Fk���;�0��ނ��ח����	 3k�w��gQ�[/Y�J%��}ݸ�N7ҺB��s�L�e���k�8��xCP��j���ش>��	,�k�#i�`b�8Jz���Ĕ�BZv%��ɱ����Kڈp�>2�̨7<��􍞫D\��X��hCU妈τ�|ꖣе�Mr�]��$��5�r��� _����`��w9���,������P�M4hRs�c�ԄYj��@������9U�TE?{W�u�B3J��o�<N���x�I����+����d�}g��X��-�R�^�eb�	�^%^,{n�6�hꑶHsP����LPN�R)�^�^\�q�u�n3-�j��&.q��RHv�K�X�e:Z&��q��S@�����l��M�� Gtw��7#
���y��_�X�֓����Q���5].�6��(I�+/�I蟡�U��48��,F31svKqrb'݀���|�11/���߳���A����k�cy:����6dJ8U��Wd��͎�A�EB�cj0'�������K��dXi;u�������)#Z�C|YbΫ�n����)����=1|�s���j}0{J������f��+^�`�g䅴X\�D@� ��L珍�R�p�J�]�n���\S�89�f�l
�](o$�Zsۻ�L�=��ek��$�X���8+3���Y	��� ���"Iq�J� �2vQ����ݨ����Y�=��~�n���H�dmNLO��Vz��dt1h9��H�V�d'=���`�K�*|�t��~��u,�	FP� �%c�[/�p	��g��9}���l<=��"�?5`V(�u;�B`1��3�3����S[�x���y��~g������҈wj�L�����: ;/G��.,�!�VN�8�������kq�"�vT^V��۪�����o�@P�U؈AC�Q���T�5p9$�z�_�Wi��#�+ǥ�s���}W�5c���@�).�i�JN�Q���,ܠȅ�T����'��p;�7��~^[�X��?��#���~�j�C�Z@�U��L��h��� -&B���#
߁O���S�CE} �6�7��ʵ�(D��<#p oѕT�#/���8'\�۠�1^�������欮 ��D�ղ�����/ii�B�%�E=���b��:Ʌ��6xMr$^.�~n+�C`����i�L�Լ�:%�^�x�A	�q��-�SZ#]M�m"��yG�SA��_��9"N
�	>�/S���m������Ǝ�vIdz��I����&[�Z�>�|=��H�,��o?ͧ���1 ��{>�̨ζ��Vy^#_�X1{T��yj+k�U�.`*���Zv�x����{�����fGM�ؿ;ڪ��b�rQ�2�Vk)>�>mY������T�+:qd��0�w1p��I]�!����(���i�S�tNv��f�O����)���Sw����ņ���1IM0%6\#[ݻ;�����#)��<m�]ͨ�³���wP^����*�.i	rys� b�xX/dӪ}�|.�ӕYg���ѡ	^DZ��Z��U�"�2�H7D�܄MV&�����L�3��9M��+����x��H'`̬���ƉcԆ�{��W��3�0���D]�4&��G�u���gS��່��0�1��9x�栌��%*�5��4X(\rv� ��(��'f�df�rG�'����8
�ӈAh���4�Q�|����3^�%bT��3!�pe�1!_�>��X�O�F����4�0�<��NrQ�AX��9BEQ0���`������Ҋ��Cvfɷ�����zr·���{��r;I�H9��#�K���4��lp�O���6�x�� ��L�h)����N���jM�l�����z�|͑-C��G>��,�����Q�D��s=r��pd"��B9��B�D�ճ[�m�D�/��F8��^��:�%!qqJc����>�nMRv�5\�#C���f�<�ٹ� �9�4i�$�1�ϫ���*��<�g��S�oPAV+��X�g���Ԧ��p��")�I�-3�i�
�8��<��7���s�u{܋������o_��}�`�_��2o��׉`�y�� �-x��J�ҩݓ�kt7М��"n����IJM�J*4�uDΪ%�{��b?((�J��G,c#y,��`YX�
6��C��CJQD��G�͘��(ܪ7)�� _іV
��V���]"�����{4���gs�)q�?�rHÁEB�l�IW�wY�A���4}�@�N�<7y����*�]�q��;ou�xg��/�y��b7�SF����~��)���� ���eӗ-)
���Vv#�q�c�$?\b�>L�#�� }<�Q�Nհ�ֶ]]ŔM�F��*"���h���"8�
��,~k*���/�����0|ޢѿ%Pe�;��[�#|�G���K����(�U�~N`��2dK}���0�&�|���oh~�����P�E��U�����B�����a��/y!�˼ſ��� �x��I�D��ZN�IR�`t�L]r�A�������֡���� ��Dtʿ�/��W?욐�Q�Bȷ�d`�|y��sNI��n �3�����thaL��Zf)����k�U��߄^� ]�9�`�V�cT�]6�nU���=�	���w&"�]��<h�����q6n�&�ޑ��jS$_i@V�D�H�����d�}���^���X�&qo�<U�v-5���#�(
Z7ý�-y:+/��_����� ��=�=�3H�߆�w�*�-A迮X�ULE���2��\���d2�������퀏��aj>�;����˽h�M\����ƅaH�&�]�-u��O��uH�����5��	�E������e�Y1v!��� ���=�o����#��,VJ�5��j��?����?݄�2�v�w׆��H������9��BVL�/U�#c}���c��[Tc ɚ�]Ũm8-D92xU9���,
���C�'7RB��>[���S�����7������?/�T&Fk���E��b�Wc_I��/*��A*l��֒c�Y�t@M���t�GG	<�~�ч�J�tQ��B�t+�dDBE��O�S���]�`�t���Y���\M��`<���!����?�aQ���(���m�5�SM)����kx�=�gt�3z�����g���Ƣk�	���*[Kk���B�p�,z�7�������o��/�FԠ6��t��u�O��JY�,�]���p�SX�X��s����Hc�	����::��z�@�;�2�$�,kuU��0�M�F�ݖ�m�%��Uq��k�-�����}6�Li��tC�~�q�a@��5�r,�T?�҆E�~(c1�k8`0\H�V�4I��{�h$��%g�hd�?�˕���3��D�g�H����
/J˴i���)�ۦ�i����%Z�]%^��/�Q�DF
S�t��o� �n�q�c'Dl��}��T!>����d�<U��H|l�Ǯ�9�[��[d���ʤ�4���O��+I�-v��lKD����%���K�ZixY_S���M�_����d t=�T�`a�v���k����2�'������� B3���&�B�gtpb�J�a%�w�kp@���i���b2xt��.l�3�xz���ߒ*P�q�gT��J`�=G>0]�����!�"̇�'b������v)N ^(�
C�����#6��A�".��%=9lx-�/j�_��eT�m��!��]���{�$Z�#�b5U}ZK�gR��ж�J��~K�Wq�D�+<��M�t���T�����k{�"�ݮ� 9�O�����}sx)B�W,�����{���oE��N�V�ղ~��'�:ɍuL�ۣ���<g��a�y�u滕r�9�#�"��d�3����'��'���XI�n$�(�򷞔�Ű��[�c��L��i7-9a���R���f*���w��:�9�h�i[� �ֲ�Z�+wu62Z}�OF&k�YDg�6��3�潊�oP��j'���}:�!z����:���SÑ���|r�0<�-����h! �v����B�~�����!"���}Q���Yxe:��`��������vb~�ND�DȾN����B�'3S-���Q���cg��Q�9���0ɹ�R��M�]�� l[��&<�w%{ ��w��R�}9F�R*�>vմk�����V���⣽Mj�לM��ŔZIֳ՞��Hh-bƈ��
%	���o9��iE7�!�ӫ�$x>ޅ��+_]T�wZR���_���[i�T�v P���ړ�c��M�ˬ���J�Śp߼+�t?�4E�F�T�4X�r�D%�4sӅ�2
�:o:T�;ZD�hF��՚ŏ!�����˶�����xAҪeP���0(NI�~����ĩK��HW����J5O>M�t�DeE����һ���&7�*��k�%���,���Ch�R�$�2s���&O��r���V���G'QG�"Q�����.k��f�a: 6��߄4��O�غ~��3�L���7�/`�ۺ�H��Bl���Ǯ���T�-���	��k��U�2��A��V�h�?��Cs(�`�lpۿKR'�/�dj�-h�=ȇ�����XE�@7�1aw�l��͝i>s�#0𑰚� ���E�p��1Fׂ��� g�Ά�EIJϼ�>�O#s���֨,m�.���ǒp��LY�	Y��������lb��]�Q���6it�83	�$�Ɖ����[���@��	��b���)�9&d��4
��lx�+ٽjח!��n�,�^����.іЛ��ȿ�$��;(����r��4Ta�/�L�r}	'=Sx}�;+e嚑-Ǎ:�����h��i r��=���5����#M�%5dc) "X}����Si����UX����>��=8����aIX�Ɋ�$֬�j��#S�9����t�U��o�BQ͹mm�?Q�xceGb��l~?�Y
�l��v05���"��ݠ7�3�y��/�[�n���y��n��
��d����� fc�{8�������|Ր���j}F�G�3m�ҙs*�z30lB�؏������P�����"8%j�f�� `v	{\�0O���G8����L|E�~��D�e�FWPJ���|<n���Z�9 ó�2����
�d��c�1~(���:㈶�ta�P����ـ$�@�&��^y#cR���R�=���0';�+	Ŵ�@�]��ꣂJ;P�Qտ; �Y��y��}��ݘK3�,�����QWH�ɋ��j�[j�E8}4ߡy.>��q���E��X7��u,�|�-�VV���z.,pp�v�����es�
R���S����̝�_@��e��m�����k�qi�O;j�l0��M���{�)�s���9Tr�?���2��H�?-��:�^��ۅ�~��x�3����% ��,����̠"����)^��PKِB�A�̷���n�Vb];�P6�w�z�[[�⺊����8]�6�ms�A�V�gZ%��Fӵ*�^3�;49���|��*y����?X�:l���g�1�HL1�~0G��lM��P��t$��R��0���5-t���Y*/�f��m�%,לm�V�k��O���P�C0��u�������}e0cҁ��$G�gC� f�;���ܟ~{A햂�O�( @uDT_�:N��.���`��𿽧�[~��}­G82�B	�k�e�����n'�C0;��4�ZOq�k��9>t��78Y:hُ��/ �:0cC�����a��B� Q��M&��{�n����.�-�y��������#֓0(���.&�2�K0H+�Yx	ʻ:d4�������f�w��Q�<����u���V��e�	�t�)H.'�o^���L���l�V�\Or��\�P���g���^�7�6���Xw���L$!�\B�Ů��k�sK�u_�m�]�n�f	޴�� �x���P�Y-�؁A$(�%li@M/�,��$5����)dj����|f6��xS�L��(�M�yT-��i��@��?�5k2��N2�E�ob�s�����}S�*Y��|ٓs��h�q�>�O��͆z5��w��(2��R8���!wW�;��C¸�X�.=�߈'�(����G/�1"�.�_�ߑ|�Gsqz��2�W����x�3B~�`6��f�/�zQc�lMW*��O"R	����?�[�p��Ek���M�`��-��{<<�o�@�(��6g����S�g��>�xq�F�3�H��3�7�#}�d��}0�2?n:w��53]ou_�@�ǜu=�"(O((���%a$�{i���} ��~,�ծ�E"#1?1G�ǚ{����#�S#f�6j�<6zh<�0�×a���˴�c�\�멂���+�&��4��а�y���.ɱ2�{][����m`�z��dũ$�4Fd��Di��f,2~!5�+�a#ɚ���O���d�C}C�'�nW5�h%CZ�$Up��\�>x� #�2��νYP�t�+�f�"Q�:�4�"=qU����&�K���Etjm�x��W<�K�!E��Ftqf�RT5��:#���l�r�[��})�|��/G���;��blH1TE;l��1�+���H4���x?����� <{6"�1��Q���@�8�ܠ_�EWA�1Ek���o�'+���v��ܲ��U+)��_�	_�ԫ�qǉ�DuA���p���TO$��,#�[2��T����-��8�ʙ|��ɓ���&bh5=�~��ԧ�� "�؅�k�6X����_w�"~��f6�?V�cB�ѕ)�T���\�/<R�(���zŪu�t�	�u_�l�)�"��ށ(��b=�щ^+ڢ����Iu�6�-��߯�hi/_,���nM4�,A�M^�B6T,�"�Î�����#E������eG�������q�U�o��5����*nd�3�TL�ioN�gl&ی������͸�q߼�<��d�u��h�����Az��ŭ_� �1�v)�Ч�����Y]��8�[�`VU�L4z2D��cDV��W>�w��h�=Ʊ�p��OH��`�U�<���k�od�͜j���еT�"�xQɌ�톹���,�W��?e��! ͅo��{=����8�9�����D9U.�x�R�>�5����v�-��Anf�uaB �Q�W�
���Y��V�I�8.����J=��ygȃ#��C�!;����Y�?���4���]�PſQ��K����bA���5e�!��uW�B�;�s�F�=��lI/Fa��sG��ī�8�5ĵ���=$*�1�h`^��:�����Ӓ�g�У/u���a��c[�-&� 豈�v�������1��q�a߀lu�[�}\��uT�����p�3K���3���WM-�.ʢi|/���\�=|%��پd�;�[ΎΑ�ҪA���t
�-���^��Z�i?N'���[l&,�w	P��AcOe����OWQ��w�;�.���P <��ϴ  z(,K�B�������T�����x������-:����>	{��$�Sڧdf�����n<��ȟ�4W�1���N���7�L�p�]�X�c�a�I�,~���`[��g¥	��aw���T�k%����gǾ�L�W���,�Ka�/���j嬪Z]�R�ᖮL/+j�]~?Z��������d�Kw�1O�,�D�G�'h�����uF�v�r���)��%d�`����,xt��BrVM`2�Y�}JΈާ�����T����|fy��Sk�A=��D�(�+xr�V^T $���&��������~U�5&j�W{�ӂ>\ϝ?˝?��ȡ�D�S��Ut#Wt9n	%� ^D��Ɠ�4���ސb�2��^��*�'Y�u�ڇ'�T��V�+��N^n�i����|��e�}#���v�ҡ�u�f�9����q62��a�s��{�l��r���g�S����
�L!<��G7�ժ���*�Μ�"t�ܾ�qf�Z���)�8B�T���L�k�!ˈ�=C�OE���ٰ����*o2��L���ķ�٤q<�,Ϳ�9�\\��$�fL��a���\k�U[RY��\���t#�pB6�m~����Y�j��G���Շ�~�o��Y�����LyL�W�(�6�}���H�#$M ��5��j�dBQ����c�Jg%WW��j�Hӑ
D��-K�Rk�\��Q�=�Cz��y4����̉���(�
0+�Jcʓ�[,�$u�-�}ƽ���o��A�B+�/F�.�wD��EE��)�ʐ�'��U}���7��i��C���4',kb��Gu3Q�5���{5?�- f:�����Jbc���ޯKM��f�C�������v�\7��hU�(!o''Wj�8.���iICc�����r���eC��/1��7Z�s8qQ���	p�̭�
���>@�հ�3/��^�Uf��X\%04
'~�n;�fNy)*�L!$k��rי��U[5��Y�o��k<̍��/�!��X�i	'�v�˝S?���>XS����7F���؅z��`��7�g
�5W�U?\�jY�d�QV%>A4�K���`#_�`� ?B�ȴ�<]���C!>����2�� l�;Q��w۳� �:	��:�Ϋ�[j��;���=�pj�#n�,�{ �y��cK��;���^�Hq�A�PuN��J�&���aCχV9+��B�h�*:�������@9���܈�qe�i�2`�1��z�����Pۣ�����#�c{Ú��R��O��uP�sŨC�h�"���L�s��!�\\����`��2j���?j΅9� ��8>[=�ǯfb�2>��σ�|P��k��Fk�L��#���ݥV2 ��	$#�>� )7�tջ�9S)WF9Q.��-~a�����+iv	�cx��Ix_�FWb���bз\��R�up��(�F�!�
����f�v�����9ʪ��
�� ��mǗ�~� �cEɘd��ۓ���.�Z�Z0ֺα'K��J��S,�9�[	Xϙ��'�@�I"qv��`R#3��ݳ�kq���U�K"8�5|Ց��[ހN���b|K�F�u�j�.9D�upi�K���B�j(|0j���u?B>��o$+I�Y�Kw�m�Ԫ����Yy���G"����B��Fv!ݿ�d>4�v}�T�����另	��aZ�I���4�魭�N��wNx�!�׭&�g' W:�f�H�.Y{�݃�ԓ0�H���a�6:2���g>g����^k�h�D�y����e�5\ˇBW���KC��t�hpr��)�ݕ(Nq�'�D$��{��?���{�T����	u8�RX���/с�8�a�&�t.�͞�ڎʠ�\��g�+>54�)�y���u�D�&��Y΂g�V)��g�l���Ą�X�s�����۫Zȳ���4M�J`��|�4����yh�sK4�$��&B��H�ԩhb[��2��4�q�=�:wj�:�a.�#6@���A&e"�So�Ay;�g4}�]J���`t�{/r��"4ٳ�pg��?C� (CUR�Q���$X��흐� �2�f����B'�'&�!'�n���qಸ�-�BfK��{�ON;��9�g�D��E��Ӝ��>�D%�<vA�Ti\�f(�(-�t��Xpd�܃�����o�ջ`X��L��i
v�#���2)�gC����8�����р��G��lEF\�u��>08oHLJ̪��?�X��C�1�y��)m��������~�+짍��v�c����T�2k��R���|��R���%F��M����=Fޏ&l�@`�0]�i��R'���/[G-�ȅ(�AO��@\P����g(����7g��p"vp�=LD���|�;��R�B�5Y�
y(���;�d�Xp5���XcX-x5��M(�����U�e9��c���I�7����G6��S������¦y =_��;���s�VU����S��=g���ȬL2�"k<�]?X�/���P�/���Q�`LZ�����r���G�*%�P)�e�,��N&<M���55��)�F�����p�$�Qj��w��i�b6b����,�c��!��'\��l�y�,�K��Ls��A�H�*��$S�q,#�\݊��{B���D�j\gt��r��6)��.�E�|z���#��Ⱦ�p�-Z>+}./R�؀��=V)�����V-�t�^/b�R0m�N��$�qf��T�&�es"��A6�\g����Gn0�r�p:����v��!*��Ȕ�c�Mhm��bsU��܋��Z��&�Q��Fk��,�����w}XB��%P(~X�y���E���S^�zrH�Q��ڀ�w0�h> ϡ���Ń;�q�p�_B����6|l^y� �u� i{����M���X�I;�>@��i;���(�������W�I�a~�x��d8)�
��1�[��H���M����\���kx߈���I� ��� $!GF��[{H��70C0=)���� �5�����,��$u�DS�KB�d-�!��׶T�n�xsX�$��<��>󥇱N2R�^�k�?#��q�w��)AP����1���͊?�4VW����妰6�5-L2<��Rt2���9��}oA��&JR��qG����e+�,�@f����L���Q��[�����'�Q�������3�1��q�UZf��\{�삿��ͅfˆ2��P^=�\B�j�^�I*�h?�e�p�L]�mf�G�dZ���
�􉾌ٺ�zl��;~q�6W�\MuM�7����4&1 o�X�9�^L"�zQ�Z9:VI��$�����p
���68�"�R]	��]��t����r�H�2�L$��4|�&h���kF�2n���
�ޞ�C�Vm��i�iR��UƮ�I����&����L�|�Q�$泉�}
{��ߋK���(Q.p���duŞ�<]-���tm�q��Ybz�'�J[�oT'3"�H4U��J� �0��(���cҩ����:Rf�"����r�&��C�p���A�f]�^f�e��I�\"ed(t���/��G�(G��迟}-sS�@��`m4�d�TJ�[kZ/ܰptg�&ٱ���������6�a�����^�D�]��X���W�Fؙ����Y���S8�2'�}Uc��Z7R�P������G[*��>�F����.���Ƈִ(�)���� ^�������_�}�ŕ*�.��@�V퓟��CD��AX��Y�˺��)�U^�t|�vh���v;\�1�����?<��y���Q�󫧽�4�� �a0|*V8=��^,k�.��?�Dql�{Y��J÷�V�cZ�"�H$aù'��4��.+���6��P*â�ψ�A���w����6(���yb�p���R�!EF+��\s}��(X���|h(u�u<���y�嫘�$R�J�"�ڜ:�Uor��tmR_���2[���c��gA�l�b�Y뷇�dyB��Ep,��VƓ3��"B�MZ];hW?S�Ȓ��/��yM�q;�ϔ|�j����3�UL���>�*�D��_$�Q%mD���WM8ݛ����A�k�	;��d�[�ތAN�FC��;�g��n��y�:\3R�s]<z��1���3�̫N}�;�z�<��d��%�������I�*�W�cn���-��&r[��s��v��˷�)펔e�7+�?�6.�9�s�h�k<�7j�K�v�'+=dfD��	]��Fo�f�-a[�:o��" C�ak�bU<¼��{qCNz��ufS<VY,���d�v@����X���@k=$�c{��_\�,/�y�g����&g��\��Y�[���Z0����)B=�i	��Eit���?������:�m���g|�ga_z���%Ҟ�w�p�~y�ߦw��n��H�k[Kbbf;��M��)9zH �Ε,��6K��J;0��Vxv
ª0\H���:A�:c�5���lg#ޤ�Ȋ���+-��ԉ��b��|�$�fniT�4��!B�HO! ?g�_�&���Լ[�Y9��e`Ɋp#o�3u��Q���0{�39�;N�E�2ʬ�'�+����ʜu���q3�����g������L�H Rn���&ǩׂÖu3�G������	qF���������K��}ĸ��+�>2A"�����T؄�A��k9W���"뭣����܆��.�"�F�mG~&�i"ZH�M?�{�|hԼփ�O}��:�.}�>R6p���k�#Z��cM�=x_T)rW����.��<��i�!s��{��sd8z��u�n��в�e�:]a� &�ZFC�.$R�%Z OBoH&:fg��R*fپ-�Z���XF����(/��!hD/���2��2=�44Ɍ�Z��y- .�"���+�~[3��ը, ����)pc%M�Ռ�b:rW/|w��-� ���ӅuJ�����З���P@�pn\&Q����*�k3[��u[�
R=A������o�alet����迼 ����8!8�X����ۚn�/t���:{Ȃ�jX����,Ħ��$��F�O)���=���	9��ϯh͓�"2CG�;��f��m��a��K���"n*h)h:���.�����ZKD�	�m�v\{`qo�?L^�	{��i����E$�	�[���U�m��W�b����,p����.tw���^�}��O�l�����k)?[)7Ĥ��u+�<���JG�+�5�=����q��c:˧F�|��fj�wF�R�:��b��������gJzz�_�xW��a����0��$}^����]��J[�7���wl
� ⢐���j�wV5`ؕ�]�Q�|J�[':�A2o����bwSc����<��>~Ձ�X׏qx&g��v����*�S?�Ч��F�W��p$`5&c����jp�-Y69���0�@β�/R/-�ޖܹ���(r����_��'�&�Oۣ��h_waN����)�����Dh�vX0��<��W���'��֢�Q\<=K�����j�G�{11�U�met�>	�xz]}g�\��mH�.����_͟R9�m����\]�H ���[y����H'��x�q���� w�EM�`+�����!ˆ`C�%��c#(����=*V�͡;gc�Bε�X*�����ΠU����axS��,-ӕ,��$����H��s�HT�� �/((��*l�R`U��"��Ɇ	9T$���F��,��_�z�*��$;K�H��J�8��v���_�'ħ���o��u��N�T=���w�!a|*�v�.w-��@V�f:82�����A~_1�������<�v��1*�K��o�8����J����lFTE�ѥYk�H{�a���v��HJvYȵ���4ҶD(ގ+� ˙);a���7X�����Q�(H�^�HU]�G��ׅ���y���_Π��!U�����Xb����ey7�A�R�T��msYI�e}�i�#�� d`��/��05�i�p��v���גf�VN��]�0�i��G_�'Pǅ=���R�I	y�Weg�4/R�\HN]#��Y�P`)d��8?q�9�3�:6�<R+�փ��7�Z��G�sY�D	�fh�p���U4��1ba�P�b���bW�إ����[�jB�h�4�����V�e�f[F�s/���i�S��6l=�c�O��$M�P+Py��w��0��&/��huxWJԮZe}L��:��5�v!�ڤRazF�p�HM6����Eo�
Џ��@� g%�gO�����	&[��r�ȗ��W�
��̨���P�rEzLB݄�"�Y)Q3�	�!!@_ roY��Z��ϊ���ʚFքP3�(��}�|���a>n.
�/��E�˚�t�W�`�o��e2�*4<��ؒ��_��ծ�Q\��: hSڠ�Гa�ȿ�(�I�����tx�'�dqɅx�6RKm�����1Uǖ�)�<�}��F�ة7�5���y�!I��|���CN:�X�v�"z�/��Q���HP�BV���E&M�x���;�Na�Dƪ�0�+���[B�F������L2�w8�Ŷ�����;"=i���ie����x�j���0���8�
 ˓���ئ͉���*U�M"P^'.��'2D�}
m=�
�Ĺ�|��/Xa�D6g]��'2R�����Z��v*�!kwYX=��>ʴ�� ԴD�,;�Ms�y�.�|��E�T�]&�fبT�|������,F�6ݞh�'��Z�Jf���U
a
K��f��ب��9]0�	95�uϨ��y�%�r\H"��صO~����	oO���"O����8�R��#��Z����㼿<�M�g?L�x���^a����:��`zxr����:�	��^��Q�Mc"|Z�/}�Q��w\q�����-����
�P<񻖜WkP� �ug��`�戶U���0�/��dҤX�#�-ӽ��V��>�p���j��}�k�K���(�F"�|�rPW\s���K�Uo�@f��@T)�!̟���	g�b��x��B<ꡆ��P{�"B�Mĥ����ɳ���K �A4���4��.������z���^6�e�ɛ�����$vPҏ���/6AZY�.��-(�F$=�+Ԟ�N��}�IU����{]�%���(|P��۳�R��c�P.R%��΍��#h��(��EA��y���<a�6��t(�}��8	Dzu���m�Qciie���4�4��0ʫL�A��i����o~�ݽ�}��ļ&��co<͝�k�Bu���C9���a���B�S��-z!�ދ�� 1X�S<�>�j#���H���n �b ��e2�h;�k{�
�7���]"��F�Y+y�A5��ߡ)1�ͭ�N_w'J,R�h@.�^�[6�,�?1���]y���6q|�%�����s����}- �i!�y���WfT?B���u*T��۸bK�>�=*���0�2�/��/����"F�cS����w�Ǟ��AS�����4 `*�%~�5f�"�خ�y��U��*d�,��mFM�@K+ݓpWZ��Yʘ�(�mit9�M���_g]�Ս�3׵�`@ug-���$@�7�� ���>�XW�c=
hm.+3�i%��yΉ�ѫ
*?6�)cS!0�pޖ���Ȇ�!���9\�.x����������Xt��~&�j!T���7�*g�fO�D��A��!��P�V�^������N:dKCb80��&d&�Řx�x�;��ۀ�LT��~=f���-�Up�"�JiwI$ڞ���t;�>{0�=a�]؃L]����甭�;�}C���v&�6ft�H#�	����������u����6�L�c��R��Y�`o���4��F��4��3&�Qx�;g��c��#2��.���	{jL�)��|G�+s{��N�6R2�j�f�8W� Y��o,�|XV�}��9���9u�s����} �2S��'htiy���e���E�R��*+���տ].)�w<2��C��h���O�������YG���rTp(�����_�D�����2?M�^_��ߩ}�ć����>8��������x�����}��v��'��Ӵ��ɧ��1���ƋR#�0�z����5	��y����`���1�;u�Л5�'?�t��?��|ڵ�Q��	�kM�?f~�FX0���rZ�ɠB��r�K�wN~��r���W�;L�b! ��~�%���z�ψ�a(��V-*z0�sI�/$��Go��W�Z%��`�
�8l)1J�� �ҩ ��>�j e����B,:�З���i�w�>�����¢I���a0@7�q	�TV3���t��AT%2I�J �-��:��T쇽���E8d[S�[m3%����)�{�w*�����Z�=ڧ�o��,S?��Zk��s��Z�$�u���eEYR��ve��� �B�m�Z������&`�ճ�Nx"�����N�d4�w��N"Ѓ��v>�T��-Up��9�"U�5���� ��m�v�X���0�Uɝ�Փ��.ؼ�&�	s)�'�i�ǁ<�$4��"ټt��T��2��^K0�)毼�8>݄��]�CC
��-,����aR\oh�_A+��kmqt�@�T|����Q����WS��Ԕ1�#z�[����v��f��-^b�䬊]���Ω��Qq��
�����UwwgɢG�:�aw��(?v���!���A	 ��Yc�@�۾d+�z<N�I-Xp|B�I%Rs�Nʵ��䩏2�qۧn �O�էS�.1����3YL��4B�DFM�qf]h@�zF�o"I�Y~/���ɫL G�~�"0?k]�=�?˕/^t[�
[�L��jJM�3��?��pNHE����?!�f&�Y�	C(�/_f7���6��c�ql,�����Ԍ�}�]9������T�6x���T|��9�n��D��+���1?�s2=Q�2��`LZGv4�K��>O�����&��]�oofV�(�&��8�i4���.I�u��űaA��z�D;.�=C5
< �m\��P�2!B�g{��
{9���ߍ�^%ԬNo�|\��Fi��@�4
��g�[�{���ni�r�$gWx��6'�aPJ��.�jP�i�!��e��M׫��+5V�U�
� {vy����l=��f9\�z���A%>).� �5��V(�	�ˮ��d��NM���8��F�_�f�)�g�bY]�H���F u��Z��2S�;�
�2��rO��×�"�2�a?RE�(�u�|l�z��#�,u&t�/�%��5��s��ˁ�Ut^���@ȍYj���8��������ͮ�4j��H�E&)�� Kx'���V�]��ӣ�0k��\��k�l*I��d�!���ȓ�RjbnA��qhFH-Am.�������H�0��(���,����AD����cI�S}
D>t�nǽ@�Կ�_����Բ�`W�6B
c	&�=��̿��+�m��1���j�>�d�ҏ#���"�:ԛ�?����% 6�F!2G��y=fhHn�����es�o
c�����`5|,'FQ�AVP��� ��*�!��s�6���0kZ�#<̕�*6IJ���ƹ��>�ez�����,�;�S-@$f�@���'��U9���B��	�C��7M���e�,U:x
�U�<O�Ӌ�x��.�Ap�7n��iWE���^��l?����C`��C^��Uf��g���آ��NC�1{Y��DD����Z.���_��^�"�3"�2�]��|!R���S��lO�����Z�z	������EC�mnu�X�Uo7b����w X�o7�s���'�	9y��:�0��A&Ʊ��te��(�峮j�A��<C ���
&�^�FS@�Cta�q��ӝ&�Ѥ)u|���^,띨�c��{U��h�I�|1b܂k`d3zǿ��|�R�ևx<��U�Z���d��#���AW������V�Hq�z����?1��A�����?����$fvS9�C� Y#�&�����~�|v|تnvE��M�3�dL^V!W�������C$P����by,i�*_��XZc^T�/�5�:ZR��V�]\U� "F��jE!������#9?��_666��j�҆z,=�)��(R���.R�T��ݣ.-J�b�N椷&�6
�8"��q�ܾL?2��+b���������#�s�L�����5���n2�){~g�rK��LF��؋Rm������,�N�Ԛ��S��*bh���,�!�C�G�;���uj�}�Ai�F����%{�@<��:D;�`�0"d�wc�cTwf�;���-l�J�V5l7��J�C$���~]����J�aY:��t����iI���fw �R�W~�l`�;W��n}[����g��%5����l|�����Z�?F���b�WƧV�u����`M��@bdc)m���7���ué��y����f�#�,p��q(k�x�*#NϹ����?��5�v�Bv��/.�:ޠ��ͫ��F�`���|Ty�ؿNxT[RKt0!ַ1p�I[����E}��0�������G-�0P����m����$�|���x?��}z�ߍƔ�^cx��)E!�Z�9�&!�<��c�s���s?kgr�v�����e��ˋG�2�o�_ݚ�l�c㝽�L�"��{��X�UЏ |Q����'}����3su�~�Z�iiD��w#�hʐ[�����4���5(��h��S��5k���%�!f�X�퓂�;�d@�����wx"��xYUݬL�W�wj>]}a�vT7T�O9%�>` �ۯ��4�����"��JV��à����\;� Y�j�J���f�q�����p��̄��ߧ�����V�8�-U��E�R�(�~�V��hy���,�b�U��L9.��b�꾀D�1��
L$q9�����~�\8V�5hR_�~>��P�Q���yQ�DIVȲ7���f�֨�("�<>�!wϛ����=z2w��L��l�iס���;,07NCc� ��}y���Nv���'#�������1b�a3��,��_�u6(tț[iT9�C;�B����{�8���D�~��P���^<<�) FjE6��TyYN��}F�2��=�)ͽ�{����}���p~��Ěkr��.4kUF����	3�|�+�Wzv��x�M�	G�W/&2.L �l����s�Gi_��d�b�V��D}=6�%�ٯ����6"T��VS��g��G�+9R�\����Q�����E/g�w��D���2"`�o��w�%H�T�0+�� [r8�p`�"'��D{}��	��=C����ܔY(;Myr��ů����Vo"Y�S!�$���0D?�O�Kp&��r��◨�'����(,|�'AkC�SzB	\����$^���_��ϕ6��`�����zq>/��h�d����/	�4`������'�7Տ��n4�9�U�600Ee�o������R��~��@������[�;���M.2���F=jĳ}?�D��#�yR"���nx0�����m1a�{Ex��?*��s�d�x��,E��Mf0^�a�n8)��wRc�*��V^�,�"�Ci�>1r�+�l�4��r?���]�T�J]v�%e�fv��K�p��5X[,��w�?�k�3��'�i��lr�2��i����\��ʈ2�HD�WcȠX��%[=�/j�.�����}�}�1b!-��l{��`ɚ��VQ�\6yII���}%�$�~�3Q�-� ��t�󡚗�Y"�<zC�e-�A���l���)��xy��fzJ�U	?��U�0)%`&���aIQ���y�NdK��(i`���a�M����������#�k51@���@{��|����Y�m�v@�ۚ�Q��z?0�Ҹ�p�O�'�\���h�@un��k6��Qy�<$��U�ۜ�[m������� �.�*>i�z�`N�Gg�E��p�"d ��?_�h��6����x�
����&��~�ˠ��F]ʱ����	�/<,onn�z�#N��1��8H(�4�Ȥ��
*)U������-}����y��k��{O��!OT׹�e^T�G�ꉯ����KFF�pA��u���_Vf��� C��=l�r
��!8��>ˠ�b�b��)z�48I]T�X�ahKn���0���2�KT4ul��e��0;σ ��}�T����	���ix^l�ؘ$�ռH�l_�l���O�|�C[�J�(��i3K��72�`�q
����@����{
WV@̜���}�B��q-�^q�r��w<�IΝX�N1<��^ܖ�A��� ��Y�������}D�wXx���%�l"����s�
YԏL�es&�5;����'�U�W9~�G��;�
�b̫n��DZ
��.���z,��:���k�ֱ��+�a�v}`��@�8t���.���J��g�xv[�	'�,r�b��6���a
��/���*,r@�÷yO�,p�G��(��~��v/(���,����oE7�]�}�CuP�i�@����M"Ɖ������`�P*+}�F.ɣ��?k_�7�rȂ��E3�.*V�r��S��D|�/,N�l0;D��Ę;���n�z)8����N�ܖ��R�����5#�����Q���@u��>�0���?tP��#3Yj�c������;�$'ǿ"�Py`�&tk���C�n�>�5�xZ�(��$����m1�DN4�{�&Ig�e�W�;�3�޼�hdb��h����y��(V��Rx��?��~V�W!��ko�ƨS�lj�G ;D`���\v����TW�k�x�%� �&�Q�5N<~��C�x����GP�Y��0���8s�0�ds�����Y���}��-�3��K �L(�=7��ݝ���n�]|q-���<����o�[�+Q[�"��g·�5��������Z������L7$���
O��nm�C��t���Z/��?'a0�@�!�z�"�C^XW��aP�ҪE�8�&!��Y�`�p���Oȵ0����m?�G��1� S�F�	���2o�۔�+�����㉘X����w�B�?M���=�<��f���F_/�Q$�&<B���2��B�
4�'�����Y^��@�5 
9_d �׊��{:��j�ޭ[���#~�!�
��e��X�lt���4�_�3@����f����x���}�IO8�j�S9@	;P�0�Sp�5ɿst*%m|\zL{���0�%\�37�V_�&��ʏ(�i� ۿԘ�sg���9J%y����b�i�=�E��N^�����a;K'{�#��3.Y���7����D�G#�b��:�.gJ�(+�����w1w�[��km��B��yi�Ԝ�d�|��]S�o"��5=��5��L�~� ����[i�����)�s�E��j3X.������(F�	߫9�~>��=�����\��3_�����g��6���CM_l�d��=�JbF�0e?�{��<vɻ�>�T�Z�CCuW����u��\�@�K�LK�ad�ڋH���^8�{)����Sw�}�E]F����΂�:?CW1Ե����5�޺�ˆ�%ƞ��-�UʟOk���V��V�r����Wl�x�����Ee�P�8���u��3m�QX���J�^Hj��O�F�+�Y����SӀ�u�%���X�x��ቫ�t�m�~=��T_	��ix|�����H7z7 ٘2  m�Ez�s��#SJ�!:V`^Ǭ�U]@"O�J[\]��r*�KIlᑚ���[=i�z�.�[�}'�I� ̺x�G|#q~7�)�a,�jVU�g��s�3ad4Y+֗ݠCa�կ���2.��%���f��ш����$��F�
l�e��)�����^%=Vl^]�L��,
A��אT�J�� Ny`c��>�औ���Ґ���6B������ʸ����R����O�~Yd,���D;���,; "}P0Dr8�$��q�+��G�e�H=<W���ۋ&Mݥg=T�����f�s\?���5ʔ8=��� 5�9}k���yL��G{nAs���E�f1��[tn�_U�*�¦���d#X	l��v HI�Y�K�F	��p��2N7_gì��T~�y�:��Ө�3</�|��4����gXV�"J�p��Om-�$c+3w����k��i'���L�c�W ɝ�¸�D������ퟓ�\�	�d��t_ʱ.y�(w�O�Aw&7�Z��@�ϡ}���Ag���ka-��NZbBA�+~�!�K��B;txz� ��ZW�BN�J�B�n�ֲ���	�w�X��&˪"��~�;x��9s��5ëb֡������f�o�r�q�eO�Hc�^vx��^�{�ie|�xKpF��QY��o4��!�T���w1!�E�8���;�����v�-02MO���ΆQ fg�?LzV�5j��D ��H�K���������Į�凯���a�%*}�,�_/n_�N���G-qۅ��~km?֎�՛V��go��C���(����0B��}"NH�@�	iۼ����5�Ia�7@W����y���@�ܼݬ�͟y��v	��^ #������g2�s)	aa,�~�2�5И_N�P^Uúm�`~>�����>�3 ��Pf�F��=�������I��rh/�������WX"wl�%�4�o�$#��H�8��*��Kxfk�m��H�+��C�+@�0_69e���'{�7\�� ��8�ԡ�$������q���ǘ�oM�f�'h�q�yFl�ƜI���)�X�}2�=�WUNy�m!ig��Ms憯�q�NF��(U�zG����j�v���g���}�[���K&��T$H��0L�8b�S�U�]�t����oY�љj�����z>�p@b�= lP"/G0-��k��\�ޒq�cЬ� 6�4���NM��WP�c�N� ���K!�L[T9+�)���k�z�#: �k���T)�M+J�TJ��A�w�Xr]]o{#��)2�-V�(|H�����_f�[�M�.�It�-��[44uE��R��(�?ڇ뻏 ,����jT��-�C�}�q�W}w������B��sy^ܖ�ͧ?Cdq#MmrD9�_��"��đ�³ݍC�`��6�+,�ߗj@Pr��t��IAE��b��MJU<������R�Զ�>j�a�����5؛ƴb�.M���(j,k�-,�ծ�,��c�� a���!�K�Z�Q��`)�6:=��\���9�Ö"]�ԝ����(��A	Ƞ�/)��y�1$N�ij{�z���n���G�]Cp -�C�a���PU,��5�b!?�Q�&O���叢�#fbۙ�kħe=�8U�i����t�w�+�����4Įqv�|��%}����C����@��~-���/�N�e�E�����2iӏ���At����"���B1.�!]����^y.^��<c��V�(~�u~|L*iS���BIx7�n�/�!��6���O�H�Թ��]���PN��u�5|����۽a�&?�@�"�i�}�͛
;p��
.����^3Dr+>��|2�������[(���9͊�;�j�zId�*�Nț�7D)��J�xМ��^]��f�._�q�1�U՗��&��5l��?��X#�����]�����H �����R���U;�t!�u�4���(n�gk�S�L�jf='����hF�P�"U�^?5MW�o���:[6��u$%����i��sq�ד��~f��R�T�����c���w���=�\긩���4)�s���u�'�+��:OBwj�-�n��$����}
��dx����{Oq�.H����D��LKRnC�a9CT�|q#j
��n��S�e��a��$V`��=]2{[w�4ы�<��M�����.��%Q��z
V&�����o�Ü�ux�(6�!���R���
,)�o��x�2��Vl��9������ �>G��2/��!<5�m���M�κ���ܵ� pؽx�t�7�ъ;����a*ơ���SS��"��AJ���7�Ν���n���j���SaL'S�I��&ΈU*��](U��lLb԰��\�0��R$ǅg{࠴W卥ĩd����C�e<U�G�y�H8��/i}�u��hIg���
)	"�5�8�7��`s�
	| P��:Ú�߷��*l�;��b��/g�0��'�a�<�ٜ������:���6w>�-� �6�
�TC�O�c�i� /F�0�^zS��^GQ6�)�����v����3�\�OhE�c~~�t�7��!)��\�7�I���Mx69�>z��������F��K�ij��R.��u�x]8T� (�q����Q�C����`�+�{�OzI�m��-p�@7C� �7�#�H��'���~
͗�~�.6#���|�l;����%�k��Vu�� � @�z����sU5M��%�J�'�NQ<���VB@�O<��3�C�t����ظ��݅��_�[�����e�O����m$�����ZҮ�n ͪS�Y1ig�k3�Q�I���Yń;��0�&�Q����%�D��Y�i��3;8L ��n(�1E��K��$�v��bN1 <�L�������_� FO�2����#�g�)H�H���]R"�7��@���'$x�;��?��U�7Ӯ� Y��"�n����ʎ�C;�|g��^�L�I�ˆ�|dm�׆�˰5��ԛg)�f��}[�o�/�+>(���$�a_��Tf�?��;>��Iiަ��j���ƨ߻o�b!���W�U��W1]��]IU���Y����xk|����~�t�"��+�Y��i6���r3�S+���yv����Z4i(f)�xO3�Z4O�����t�y�hF[)���Wm�͝L���s��3^M�P)��2��4��/H��×P��ս�b�u���Y�q�{{7-��u�جu�3�s�TE��+W$?�NX��ʺ�R�xb�������K��tH�ԣ?U��4�MW7Ȟ̨��S�s����s� H��N��$/bm�5�?�X��@z	s�p�����L&��Ãb����КTe�r�)���s��A[2c�0;�[� ����s��h��5�m�QN�����t�y~��V�Mj�]k��̄�<�!QDS ����(/ԁkhq6��~����h�X{>�N���9�1rB�w�TL��e�. S*N�_ސ�vW�oUH�y�m|�A�t��,��-����^
e�\�Q����:�DG�����
̶$�&Sxh���:y������2)/�>�A�P����y^:�~������̾�|S�1p-��3�1�E�))�D�K!`Q���3hٛ��8i�!B}�!%(�_i�Ѝ��p�FY��8ׯ1H��ݜr��߬E�l����3�fg�!&Z*?A�D�����]IЛ3��$)Ⱦ�n �����(���H+�I����٭\�:��� �c��$I�G���B(��>!}��P��{�{��s�D)��\\�#&]Q�>����|jƱ�8	���3�FoX�)��k��Ꞅj�j�N��lߟ_-���4�t.hl��u� ��:k����S¦0O�n��͍�"'���mZ�jMy�����ܔ��BW�"��G n�+.�g�r��d��H��I[x�D���W�H �n�$���-=]'�#07N��;� 
���E��C`(#!�J��
5rb�s.��8�FW��"`����[��CU�8�G?0A�l��������	] ��o�NQ�tx��^�&��=�Ĉ�g�/1�p�m63�&�����	+&:������p��x'İ�:a�B�U�i����gI�mdBB�i[W8��YFu�X��/���=��ĬMw+��s�fOQJQ�{M�}�lg���C+�W&klfwjV<��{�/HC���G�E-^_R���ҵ��EE�ml��,M�<t ����H>&�3�g�-k���X&ѧ�#r�^o���##�t�WmE�e[b�^���%���p��퍈j�/���&�o��u���mC�R��K�P�+x���D!D�('���X�N�X�O���%�bހ����ɨ.�(�Z�F��jg�Q*2]�e�����P3�v���A����Xvi����b�c)��7�}|d�DVAV�r��`�Y��;I�m2uR�̆�,e�Ɉ2&���ê��.��!Z�ͪ�?�Cҩ�0nuH�|?�i���d-X鹣��|3M�1��b�*�e�y����F�	�[6;���6y�k�"�f���/u%��Q=y�����[S�|NC+Ƃ�[`e4��y���kl�&� �|����!� �����vb���=ŵ�ɹψYDײGX����&T�>Jt�"��s����<�E2kg��z���'D�!kQT�HD��%��/�7��B>k6�ԪTf$R,z��a1''Q�kH>��˶�}ZAW`��\����L���� ���&��/���#���	0���˫��N�@���Y��}?f2p�h�W+\o���K�
�^��Y:H���N� �y"�ZGJ�P
<�~��.E�z��2�sh�Z
�����g��	��c1������pOO<p(	�R�F�>���m��Z�U��*��o>��遌�����|y!�O�&�A�a�D\�G`�li�;�4�0�!桡꾗�+R���W��� Z�)!���={��A��ì��"�	X��Hf�t�Y\�`&Ԥ��KF��!���D�����O���M��P��R�_�EA������xb�-w�ӷ�~a��(;z��#�Av N��F-1��P�߾2)�iGw	��2FO�IE|B_\�!��
}t�x}n��RS�t.u�>�Φ��1T��I��H"�Qo�����W����&����H��q �x�v���7T�6.�V�d嵐P�����7��e��sU��~/��|���un(��S�JEݚ�4�cv��Q���c���u�W/e�V`�T)���t�!z`�]
.�_lr�Z��\l��P�Iv=!����ٸz�=�(q�����8��w���G+z��Nw#��pƹ������?NH�Ïm ɢD"�:�r���ʞ~��;飡x��Eli���j�;�R���=�)�.����X�(y���G��=�w�|��pN��E�(��;_���4����د���R��[�KY��D��B,,3l���;���;�]����;�J%��@^�KߦXBj����е������O#��[�Z���MH�Y�
 ���?D��yͯD	iF����
���UҠ��闤p�A�C$k>�t<r�Y�mG���qf,A흴W'��~�%``Eù$���m��qjr��7g���16����:h��ƻ2NsW�Q�AU*4ɇ �0�Ƀ%���\5����Iׯ(c�QRs����˼�]�5�Bu���x��<0�{��I��WX
�+�����BY�^�X/|m���84�ؑ9�	s�F=���ۑ�d$����1��
[�3@M�{���:A&|j<�.b�e�c��}���2��Z������<��VW��N5�\=�+L2���I�i���S|۶ Ҕ �O)��j�A�u��10�eW�^I�@�u���L�W!4)!J��=Gc�˖�a��b������!ɟC�!�QF3"O���8ZyA�y���fm�M�#�c�{h��?<� ��E8�ޯ������-բ7lq�~� E��J�1٬M8�Z�j�t^������M�����v�R��]lg�f�vo���l5w#��.�Q��/y��&G��"P2�h��ڗ��_O�_:��6b������G�c2KF�E�1P;_U�?���[a�w���3K��R���H�cՄ��ƉN\ٸ�W|��Ǘ�=:�z��e�,{J���$F�>��G� ..)�ܹ��l�16�e6T�'?�)����{�7 �~���x��� �
fHJvh&�T(�q�:p��u7en�ۙ��m�D#�8��N=�w� E���=4śM,zH1Nr�7�H��3 �Nlq
�^*=���E[ޙO�r�JKV촪�@��>���(���Daj42�$�=Q���!��������H2f�}1��X�k�m�I�}aݕ�R�4.ֿLE�^h�d�WԂ.	�i�*r���:h�e��������������(<0�����v��4��g��`��'�ۚ4u`��t�0S���-p�|d�8)��NWhd��͗���H	�@�����Bf�/��ȹQ>&�d ����,���0�L�"�+�"��w��Ri?Fgg4}[��)�����#�ũ�0���GbT�2��
Z�8q�S^g���]�������y��4\N�)�P�m�%�:!�Q�k���+��`~X4���H�� ���:��X%푛�Գ¢�cA/�]�L�<\jDa�X�9K� �b49�X)�X����2��_fW�j,S/:OZ�鿜v�^�t8��#ϻt��dV9���/�%�#g~�Ny��F� �ib�P��Qt髨r<�S�!�ma�y�~�Mʾ͒@��4��;f|H+��*@i6���vH�B��6�QW1盃&(y54k�Ү��Z�F�Ě����/��~~����yc{h�"�Ô0s@��v�(��v�{��
�xZ�pэRQ��M��"@��`,'��&��nΗ��_ħ-�2C�6��A:���$�����j��F�%�}�D�R���>�\�'ͦiz�w� �-��zL�*��b�ۣ���LKW��A-3u3#k�KmTU�;��b!?�t���il�3fE���S~��t��FI�f�V���1�mAs+�U���C��[3��+>�Z��j����w���N{8rD�U��=(��w$�"k_:���'؀K�%b�1Q�*Ut?���h��s��]	,�HZ��x�_���j&߈��[.� 5��I������3u|�&B,+'�z+��i�*}��'�ݼK�xB�F��,�����f���q�4�?�&*x]ru��E�ɐ��:���a������^�^1����q@p/�[�Չ�`����z4��Pr=��3j�(��V�z���GiO��A��"��3z�
@�TM>-|�.�a��S^2q�iQ�$�l����l�,]�A3���E���2cq�B�(ޝ�,�^bU�í�����K3�M�\��o�޺�=��G
Ֆ�P��Ō��MxV��m\Es����՜�o�$��8������owmV�/e�i���I�飖��8\���Z��]�D��8�L�lW)'��gB��n]ɿ�����sm弽"6ip[��{U>&V)�z�F?�o�g�N���&Lō+��,��=V<��N��Z�`F4`7�cj%�	�7����w������V'G[֢P��yM����o[��rG��N�=D�R.�~�~G��)�"l�1H�<���K��W�?����<����y���P6~�:K0��,�bI�� jy��"�r�遬G1|�N�dG��r���|q�Mw�:�.g�FA,T�p��y�s�C��K&�s%\y���_�����SBA�)�����_J�~�Q4�*g4߳MF=z��0��ݓ���砿�7_��ߏ�a�#�w&�B��ψ�Sa�,Ew��9.|�bN��<r�]����������x���L�9+.�J�Kf60`�T/k����t�-?��A�iI#�c*P�]�Y�E��없�����SƆ)/���E�� [�����"sr�����^������3���neJ6�Sv��A����������Ϸ���*�/�W+G����36���cP/�0o�I{K����I���U�����曂�aX*�`v�6�r-�Fr�S�A�Лa����	i�|�4 j��/تN����6L�1SV�/g�+R!&��m��iEݠ쳙nW)�#x��m�����x�����Vϐ]����������)ϫ�V����*�i��3�����V"�G����K,����U���}�����Q�_:����=���P���4y2H1�5.���9!��[�x({�	ʌ\���_�-g�[ⱬ�e9�J$<��2�Y7D�=��8�8��y�MB�y����� ����ϊ��
 յxL�2+���U�w�� ���B� Q~��pz�\�.9@�4�������;-X�!��I,�W�c߾�b1c'up;��$J O���|��8dR��@dv�͹z�k���8zT���%0��y�o�|�S9�A45V�Z{mH��v��͔e&�.�}��v�m]J�h`?_;1jr!l؍@���W��o�W����f��ہ#a.��;�5����;�O��E�9NԴ��5ObE�D<�s	����NM����)��tN�k�� ��(�����yꜸ��ܙ����C��ť�܁�@�JH�:�������k��@i�Y�}#�=�Oc{��zRb�"ܬI�9��zbN8�=,F��9�f�e�z�B�>��i�?Ru7�i�)�^J��N��<*�%�����H�`m.]g:��&�k@�����RR��?U���n�e��c3~^��D�U�>��Q1�GO@��.��p7>F��7��0�r��O,4�d}�_8�m�+[�իޏ'D��F��M�*� :<��7w����ߌ˰<�t��=Wn��� i�����/I<a�;�봑�ڽ��6���%��G{�SW�`��L+N�Dc�����ýAP�IΠb�ɀ�݂�	�ieuי��u�l��ɪ�7ɒT˻Z,R���S���/A|��)�޿�� �7�������G�m;2`I�Ϳa�ѬT31a��[�F5ʍs��kk��\���pe��:�U�/�R�K�5v������P0��y��C>�5S��y������b3N��\��/:2W!��{���k0�a�#\u���4K��4��3�(=7�S�����3�MR2=�d�hO$�L��!�x!L�X�Խ��،�Z��:�(i�,1���<�s!���0tМ#��i���<�7,�}$�ҹ�K�Do؍|��ml[�R��j�dv�p�u���NK�c��$�n65�!c�M)�����d,���x�6������u��9C���!)=��}\cPC.��}��E��k�i�!��2�Z�1 N`�<�͔�ʅ�$��W����Tc�w�fځnN|Xj���2���4�:�$�����T�%�La���{�8���/N�$��XmZ�T&��oI�l�<X���Q�}����ۡ
�	��·X�ٮ�d�星�֍+�0~_��	~�G��itU�A�Hi��W�lO�a�մ��RUq4xƓ�� z]�|�����昰�2
��7i[8
���M*9K[@�3�M.��##@赬��n&<w�qt
�n#SzxD���yO=�իW�(0�D�xg���!L�+�������[�j<��e�����'���z�O��Kˈ\vG\��z�VpE����x�"0f ��Ըj������eë8#��=K�����J��v>��
?�(�y��?�ete*��K<���V:fl;O:U8mW!p�]:%�"��gG濇6s��TH�N����y�� =�нLq�st��m�3���#ck�M�ĝ2]R�'�&鋔G��͆29!(Gv�u�%�v����/QI㿟�P��HA��ˋ(�ߣ�V��yf��Ӧ���v&��	�oNt�dJjI4��4^���3\H܄����B}�l�AX������5�	v�y���>���M�I��`�C���\ދ��_���@'����[Η�L���ʊ��g0�m��@` %Dj�[?:U(��M�8qM�ſ�N���f=IK �tbn�G\��-��Z�k[�^8��%:'v�m|��]"F��"��oh��"�y.KdHV�	����!ù?8�d% ������rb��痟�k�J�B��'�b�CLxAD ��b*�������J7�_5��k���o"R+�uH]�`O<�~ ��4���jI��ۈ>�w��F&�p�N}�<�k�ߣ�(SF�e}#���Bb'aCִ��Ц��`>^$y:�j��M}Ӭ[�m�H�s�p�?�n�@K�u�[DIhg�N����s��8������K�=/̖9�*��|�ޛ�wP!�ʭv�3�Jdd�r	㩖�3�eG�Z�Qv5ꙩ�o~�S�����.Ӎ�'@<��{N�R	?�c�F�	Lz� ��3�R����!2��Gg��sJ�n�(`��ߏ�T$���t�`6d:0�����C��$Ǥ)������k�
��*�#�Y��&�y�gr�	IAl�6��������a�c`¼z��T�e���Z���v��؜9�k��e�>W��Li��^}	�� ��D�y/����,Ab�Vn���Џ�h]�M�-8�d�`�N���ƚ�ݿ�<��q�����ϑ���ztxc��Fm�A�P奔$�PM�(I�Sh���ٌg��>�i+Z�����PIڼ�j�j����Z�O���5�G6G�\�P鵱$j�BO�$=5yZ�ZM���cb�*�d��+q���Z��RT9V�1Ac��ûB�EBo'�-D��q���î�%�Z�!��׳�m�rB�m�7.y��is��? �IUsORO���we�����3\��K�߆Z�y�-�Ph ���p���`>�J	��bv�� �ǃ�=�ُ��m����1��"��-��j�W9�"2����h��1ΰ��-�����7���DVՌ���x�rS�ƫ�^�"S�c@(��0,�1� �<�@JH|qh!�%?H{O��ly���A�NXǱA���'�ե><�>������#����RX��@��ᘺ���§���I=�%r`�T����,�[8����s�����(�J���-)�%���+P{ԙ%�<ʬ*����YA/ĭ5q	�׸п�R�h�m��Y	�>&ŗ��o�F�d�L�H��`:X�z��U�(\�)�ɷ����v�iĜ�/70������w��wqq�z������E�yvT`'���b>���^������tS�+�1��A1$`ӈJ@H�����,�������dǏ��;�:�L�NI���%5�覞�G M��f�*o���t>��D����\^k"��w)�vA{lS%p�-��j�i>�g:ˆ�7�5�gߘ�=�$q}u�eC.��fׇ�^<	�Ŗ�d#	g�w�;S�L�%}���CF�4����)��V���YӖ�[<2�EN'/�f`���ihE��z����{��ɈC]e�����0'��E��=*E����h���IC� ,Y��q��h��J�᎝����j��7�3eP��_cӡ��^�!�� &�F?���I��%c�a�L��>�,��ve�\�tSt�~����eY��m�w�A͐&:q�p�8�ɹf�(m�bNz�ܱ���~�؂�8;��*��&̤�\4�Y����j�@��\��B1�u"�j9���^2>���9
��T��$v����(GQ�
�ö���F�Rb�����0F��}w���/�Z����U����=d����*��[��$���w@�ʹ�U�\��/�Țh�U�fm�k�y�%����q"hUdxo�WY�&�6X�j�����wA�k-4�
eF�;�iO�NDYùv����+|sM�DJ�q� 6v�fb�[֨;��>�t��D��_ؿ.�z��Q������J-.Z���!T�'��8@��pp	�x�س����u�����;�ϣ�埢'��g�����{�����!�꽠Z�,\D2�2��2sLR��hv��)r��p_5o_�=�%�)����m�����[�s,��Έ �^�aV[���R(��`���sU��|Cw��l2�B�dk�E�2d&����`HV<�Sڹt���'c�jJ"ALQ<����Z�� y�\�Eu��H���x�T��A�jX�x�f��a	Lbx��W�<��E~zވ|��߃��`�W���ݟ"�=��/���>�OET�@Ƴ��"f&���g����I�ۊF��~~	���ǵ8���w\�T�,XZ:��l��R��5D��+u�s��[���%f�}�_�s�?�k�I�,����6��tO8�Y68ݜt��7R�~�a3S)_�+L:���	Z7��d1������B��3�E��Å6#���q�f�12ėiY�ϣNko�~�Tw�b�zeG�0� Ä;5�D���Ŀ'U���t�#)IN�q�W�&S�6�`q,ݑU�'0QGv���M}���j(r�ʺf���y�;�2������Y_&��SZ�,�Ϊ�XQ�ѽ���Ƚ�r@��Zϩ8k�j����W*��4�cug)th�ۗ�E���|���:'`�1�bE{����A�UϺ�Exi�KK��� ��D}Ty�Qx٬;��T��:3�e�#6Bu�1,��]GqL�����,��B�����1��9���syn��&�jW	,2^l*!ī֊v�u�@$��L��(L�[����?ooE#���S�E.x��:-��l��-����7�I��9�j紸��vX0�?����n	���&p���r�F�k�!-LOo@�|�<p�"|Y��QK(ڿ�!�3�6Œ")�� >�<�Ǟ�J���W�-9O7�WQ�1�#���n�s� �+,��]�b�M���EH����ALr��3	�p��S��7���[��=!öJ%����}�Ѵ|��FX�0�����NbDo�dp7���`�c3G�㽐��S%����U�d c��������AD�j&�U��=U�/�w�++�B�#�!�����4�k4�tcÇ�-�����5���O^�%�#J3����w�V����;�0�s�r~�^�e[e�e��Sc/y�����j�XZi�/�8}�+B~��2t�x�c@$r�;���m���F�i�B�%>��u�.�e�<@� ǅ쐨����ͼ���i�|�?*Tu<���Aj���K�b! T�Ww򮓼w���8~��Mq�	����C�/nj[�,ܔw������s�Dh�O�`�rU���jC43�������Q�uo]鉖i�~����	�y��O,g���e����$'��I�.��D�G�/�b>}�?�z�IJ7W�h�F(�X�X��X�RN�xH�t}KXݲ�� 9�V���̊Hs�c+ �p�"gC�od��j��i��%���H=�7�x`-�I+�GZ??ׇ���- �����v��sx0:�����ǯ�����W�5���� a��BS�������:�,b0�j��pԵe���)#�,	�����S���YȨ�	W"r!/ju�6��5��)����ЯS�2�Ý����)?�b��K¼��q������j2|�.+2��S�6YT�����O5	��h	Զ��"�y���\�\�T��{�9J�G>�Q&��'�!���������A��w��ƨ`ڡ�a��ʗ���G��qn�	zx�e�[��W;DMI�!-l<FRBl���;� �\��O���U��g�p�GJ_X�%6$���V��������@��H�w뭶���""�H��P7�HܴC?~ xm򣚰7żOPM�l�I�f�vL�YC��i�����%�RcMn�C@	8�J�����R6,���i�F�Q�|���ɱ��d��@���Ȣ��-���0���������䀸Iˮ9b�� Wز�=��&Zy���߾hm.a�d��]��mGS=/��Q��<�i�B�UkN�S�r�&�o[Qz��z�a�C��D��E*G�I���~�|o!X��^-Di��y\�D\v�:��tz�N�:6�0��Ε��E5�m7�)�>�r�Ops�/̾�x����mR4��y�+�J|k�𖤥�<v�*��/xFtN�]N�\�-�����������O�JN���J6MΊ)�(�w$�
�6�	��~d)jgy�@��C9Ye�Q�TM`�1Aޓ�.��;Q��x۲y��w�������ո�X��^�������v}�34���,b�r��$�n�^Ƹ��}����r�Z8��]Tb(a��>�f}%0�.}����ԷA1�`a��c�.?��t��fD�Œ��T�Z'!d\d~5]�ڕ/���F����Q�[�U�gz;��9�ޤzu)��s���~�b9������
V`��?�B��3�k�fg�mr��4���x�9�7N��ٲOշ�#a��zNx.PW����(+`�c+��RZ]E$^-���u~�;�����zw~ M��mN�y'q.�,갢v�+*+�fmU���o�U2��В���kCuu�9���ı0J�!O]T����2�{�S+f��{�}��7���#GL��uh$G��I�B����vEk�\ozNY�V*`�V#�wY|>��
+��LxI����8��V�R�N|
tui�`���@�A`v�̫hE��L'��1�K#�A��� 0 Q��geX6��w�[�v�lV�ҁ���H6�-f�q8߻��B	�� H��[6�B���r�z��[L\&S�M}`:�e�1�үw	H��K�N��!C�1 Z����WB��Ҋ!�oӪ�4��z��VH�d]�dy*�_��p�	>P��9�*Oj�ʢd��_�=ɋ�%�Eu�K4��}�a�-PZ�G ���R���<I" )n5�qv�J�Z�}ok��oZ�cM����H3J<�dkפ�N!}�ݣo1d�z�ل�dPjJO�wouT�D$X�rLOW�j�,	�!����R�0P#IK�����;=v��j(�b��z["v���V�<#~�fD�Q�TM�1@ ,Qybӥ㱣�0+�MO�	�)]˼��KqÈ��.x$�
B�>�Q�S�p�Qr�������� �B�A�u�D\�y*Y��S�w}�gl*�<�yB�	��!Gw��c�s�`��l�K��3�Ow�9�	E8w�2j�Re,^��,�H+��_�ab���%sY��ғ��H���U�/ʸ��#���� 8YƋD]��t*=D���Q���-��T�cU�G�m)9i��\Cݬ�MQƳ��'3�4�E_� ���rRs�ss������O��9Q��9��l�S|���a�"4����D�JpU�wΈj^S3�?EqD���kER����h��d�c)K5g&��%Sj��?T`���q�?՛R�*@���e�>�V����9O.-Ah�##���ھC�M��G��_�\�K��F6����2ũd*NE�XL��� g��8u�c�<���=ܸ���|x�o,#��#f�	kw��Y�I�׃� �'���m4&K��ag�8;vv��i�2)���|���F{���\%���/A����2�ヰ�:����=,����(�]�V	W������y8�3��򂵕ˍ�۠�K��@�L�K�R�(G�Ol�����fơ�h���9Y(��D]�Ԝy�!�e�	nD�7���1����8sꥣh�LU�! n�ͷJ�P>�?���I��6��5q���u��ݾB+������WUF�~��Ny���NͱC��nԵp�pKU��dHLwyD�ͿA���:���E��P�O`u�C��c�e��2=�C&kr���G�~�~9gתCaJ`)�gq��vU'�����I!�&�F��_y����Hzxa�Q�&�lž� ��Fݒ�u#�q
���t2ȉO(^pԙ�n��D7X���|�3{�΍�ύV�Rf]-�E��,�]9U�!E�s,h���kT�L���j�j�����_����qʼ?�("/p�݁/K���������y	+�j�܋��cHr<����)v��ŉ{!�Ol�s&�5@���AQ�޸�ρ���ܵ��:7=!�8�n	�}�{w7f'��c|��%���Dx]w��C��K��}�V�h���,bZ�2x8�QN���I���OOi��''�M�/!�b:�P�;GJ���83�j��c�&X�҈��-å`?䆊_������ݏe��G��jo�.�]O����e��s3�@+�3+��˹e���w"�$����4��`��tT&&U6�^�|����C�'�4b;4R!wn��3�����vsI��͜�o��Ms3Cd5�`��@����X���P����s��7��4.$��'�Vo��դ4�pm�iW�e�"�G�!]��Eh�Ƴu�%`d�|��7��D"D@8�Q�*gm%b�.��|�uf(�&�T{��x���)�=)�|u_ml��D�]��K���7:�n�5í��N�' �xYUc��&)a��9��|a/���ۨV��'�lJ�+�����3��X'n����&�1 h;S���a�����Bs<�'�_�����"ͨ�rԉ�
m�ڌW�(�S�ׇ5h�;�_z6� ,�@�Ϲ!E����v�8��B�����6R�7��Y&��\x�����T&������I��н�H\¹W� ��t[u�Y��o�^�4y�Fr�v��Ɨ�^��]=�C��fAj��4����:R�i���F�O�h����+fl�:Z`W)\7�I�C��6ĥ%VL�g���x�`���50� aԣ�B�O
��+��~�)<3��o3JT�h�b�.�܀���D����q�����,m+��h��@���.�'f� W���%�����"/nF"4�R�ew�a<.>x߹�~�|2�Ye���`))�"��V�!���5�=��s�O�PE
=����ݓ4�!�yk
�rD�(?��$͹�΅abTBb�P���`E�O��q���=;1�&�%����O��w9	�o�P��m�A����7"u.��ޕ�Z�raQ�F׿��l�0QA�+�:�85b��<M	NF���!�QJ3�vy���B㶿��ܨ*�	 �
6�]B�S�o� ��2�����1V�J�̱��m/����dduۻ� �>�
"�Š;��|����AL��I'��"�3a@#�?�M���ӌ@�9���s60��,�׌~��ߨ��sR�A�XM��\J����<:Y,�C��\@͆y�~dC}�:������8��{9�ᖠ���B�Z^	0�U^��c�^��T�oƵD]H]�HF^<{dè��O
�� !�� �aO0�h�nv����J�Х�jΤ��!���1�ҀKΧ:A������1.�֖�z����c������Y<�W�il�p,vb�v�FM��b� �պۯB)����8q�V�?J��|�^t��4��r�����ʏc�ѩ�߯�
�:�hN���c��H&��s��9V��:�����͕��,����$Cנ�{���Յv�8�'Ʉ��8��9�A��!r2V������'�ȍ3R♏���[�[Փ��&��A����rh��xűyr[��k�j�g���~ʍHՃ^w��3�����.���l<,������,����r:ߥ�oS�@��agD���p�禍2.*E��'�X�_���W��$�Q=a��,���an�[�v��HZ�d�K��.�s+Ke\��y�^+�I��*�֛hu!P��\"f���dn���VƤ��!Y;�遑TE���e9��i���8�j8y}Ʀ���X;���\�7DM ��o0@$ue�|��;]f����.n���R+�=����\��X߃���Ple��F�7��8_5����`���3�M��(���x���L0����5Pi�Y��"Yf;찚^���h��_��G����YS^�1�7�Cq'�te�H�ؗ�&*���5���/�S:b���_�\��d�q�k��J�H����6��kd���d���< ��\��ӲYf��fG[h7�=�/M'e�|��[�f�I$f';�+c�w�HR�ݎ�;bxVO���[��[u7M!�ы$����q�XL�T	p��HLq����|i#*�U�[�tP`u�tg�H���M��#J�`�>a�l2�2�MZ�A�GiXs�̗E�vh��?�'I$���a�������
�̱K7�ܶ�S��e��)�?���/=�T�Sg�+@����vāC��5Z'%��x��f���H�\H��;"�$���KC!�������sHg��It.xka�L�_#���o�Jп31� �f6R{I��Q"q�[���t�Qj�1�7S	�]_�'�ZRc�b��zL���)��]E��^�Q[��2x@�o�"Eiy�(��>��{�?�U�"f�_&$�]�&H\>w�;��|���ͷ����Qf3uS��F���X��# ���哙>��2va��T��5�B�8r�ewq~�/!%��ԙ���h�G�_;�{TZo�H4tH���z��	�g2��h��r����!�b?ya³$wiC@�,&���)53���w -�DSu`�������^��YM���^P�I�$�$OOuO'O�H�u��]���\����={=��V���YÝ}(��#�b$���*�J�2�bȰc|"�/�����&����1�o,�_`���F5I�X�@dW��;>��9'���6R�AG+�$4�'�����TSDS��ɝ_��x�=��ب��|�]�VHa���������$5oGT��0��U�w������I�r"@v�T~bin�	�}���Zl�r���>��e ��}�Ul��=���MxK��<�6t��Kިe�I*��j����ox�������5���RTsL2e�9��e)fʯ�Ȼ��C�}�_�9�z�������;������)�j���Fl���'�P4�o=��Ù����V�4�Z�<�kzD��ǳ7�7g��ɳ�!&�@�
߼��=��{�0�8��
�q�u-��Ĭr m�$��_x陌<��R^;+�=��N�ܖ��I��W������k���n��%*��m-9	��#T��()q.q���FqT{ ��i��83�Jm��dz��t)�����7ܧV�A��X8���uf-Ҕ)��qF۞��F�q���k� Ar=&^�,q���,��q-���GS&�G	�PeƸ���*fl��N^]�HD7-P�=b҃9ZK<tx��>j1�1�|p���t��ON_!i,�9gd/7������;�-X�B�w(, n�b��zU~���D&�Bn	M�mp�������|Y��m�1p����ͩ(�R�h.Dy?k &p�x6����䠽��yd�� 1�}5N�ki7#&]Ә�_]��p,|z�2�%<�Q���T�Ǩ����2s%l��EI����Na�X��5��E�{/րV\�8b����%l�+�%�������s�(~8f`%ݔ��RQ�n�~l�����,�{~���\�J'���]�FcU����h�=��~]���z#�
缂�C�!��0�
�Џi�n����� �i��o�C��	�g�I��9q�̮._2�{�� *��Wa����L��[�֨=�9���Ǳ6zhP-��7���^9A���K�x�~��`���Ɨ��j�g� +W�u�h�S�;Q=L.��t3����h�zAi�qrAR�$%b���#^��_K���1��r�2`��Ǎ�ڲ�A˴�.f�}�xE �l�hc|AS�Aĺ
���_����+��_'�b��)�#���,���ȞcYb������l�����3�0���?p�'*�~;f�d�l���dK�hed��f���R�Y4��U_�6��t�����!��ű�·ܘ�]���6?`�����r&j����j��st���V�#�Ԥ�}>7K�v�It�Ϟ�(-v�K�e*=�oD�=!Q7�eT��g���'7���Xe��
��C�n��m��>����eJTd/���@ ���t�/ ~���-�D����r�x�>����n�;�pDcFe����n9R'#M߂z���'9? =���>�{H�oAED2��/d�5�]�&���b^�x� ���d��O�88C˛g)����"����k�Z��n����V!��+�2��w��@^�܍ G��x��#���E��d�t1�t"�mu�$Ř*�Ⱦ1�n�m�^�dE���CV��o��{� �I�v���
���=vj��`ΗP�e$��ux K�0�o�.���ia���9��3�JB0,�P���H���@tbQɈ�U1ľ�:�ِ��B	@ݢ�����T���h=� �턁m�;��V�y7<.�߈�T�74��[��s�r��R�8?њ�3�xu�2�e�"�0�.�h�B 4V�G���H�!Y�,%w_ƐTNϞ���Ee��\��sc�l��iK	:.Fo��$�b��aZ�K$��|���޺��F�r�(Gp�T�x�!�t��I�ݴ>��E)��6������j��ֺ��=Ze�Q����ޛl��
ƆYx;�?��]5���e<Rp}�M��Q�k�LƸFf����|2_��F%M���a��Oဨ��=%Tw�;`jlX�7I<8��QZ�1c���m�$��b���'���Q��y^p��f��L�	}J�#C��'"{�?ТKG��͕cnM��`{-\bF�O������*f��큐���݀�����
a$)�YcT�?�m�hH�
h:F���5�"����_a�|Դ;�w�;�ŇKW��Z͠�Uu���s���� G
?KTyM��K��6�Zj��Mˀ�hͬ�-�d$��J&%y��I�hQ2�V�?�5+3�i�gQqF֖^�k�B����9�@xI�f�)�*#�C�B�T�dS�q�dj,Vu'Gz��qPyK{�/`�Pz�K�^	>&�_l��/|Toy
�Lm�a"�9L/g2�"�H�kZ� ���ˊw���n�h�
�HJ5{r/f�-)ns�ځ��nr�s0=��,DQ�C;���8c���m�󌬾
^1ߏ�3cMb���o�b�-��ԓ�
?���D�7�w$ Ry�v���Gl/�9���YW��T�e�0�R4r����&z&��V��$��쿾��l\訳6�(��Qo���h���l[)�����1�땵n�`w|&�W l!Ws��I�m�ؖ+D��6�°e�I�QЂ�`�>S )�v'�43��U9qeG>�7XW�8�?�Qr���W�F"�a�qi��zp�sa��ʆ5� \Y�'�,��o��4�=ዯ���k����H���5��4_A����}��9n�E��li�
�v	Uf�(����Ɂ��])��T1%�+A*�&��M-��
���V��:f�T�`a9�n����S����g���==����	��˽F�_�>�e`,�_��d�)$9���s�/�ʕ��� ����-�? q�T_�
�݅�@�Dm��;׭3%�=j��]���;�4ɤҿ�N%�����ٗVR��Q�sF�'����[���Q����<��}��ۉGe�S� �`��}��O-�2RX�Y��ʾ�G�8!��]
Ћp-��e}DW����e#&��l���΄a�ej�b���؏r�͇D����p���g����>�GnR�P�R����>�u�xm)D���b�X{d*t�[�t9����s��S8��'�a�����88��e�2[Gۂj�\�4!�UT�q`�Q	���"";/��pDEz,�� ��쫱�T�݉*����zp�ƅY�������N��C���\R��V�Ke~�s^���Ȅ	�ׂ��{�~���n��Ӣ��.ʽi�n��?0�yw�,|�����
@ߣм��#k�: ����^�V�rK��(��s�7���!Z����V��&��b0o�Q#v-ɕo6+W2��X�>Xw�C�[j�j5Y�Q2��"�K�dd�)/����Z~������2��~�U��b�B��1��s��c���69e�}1�C�����<W��Qu��ݕm.?�~�x�
p��2֬3؉L�&��a�/.F$�Wb<(ć��h��o���|�cGD�*��NЩ����O�(�7L g�r��V� �	������|��&�i����s����x֓oA�u��!��^kYk�j'�i߫�F�����V��Xv�2��NVC��x|[-W�o���N^+uK2���[��S�Z&m'^�pʖ�mm���`�����A�տ5k�N�z�.z�=WM9��1C~H1�TO���v��*`k��m��(T�g�I�ѝ��9��a._��+�x��Ӈ��XFϻ�t^\���Yn%�!r�L�{.���"[�i�`w�:����}��C)����	 
k���YNr���|(��I�����0�J���H���x��?�vig��NP&o�~^/���]�>�f���F@��h�+W��3��V @�M�� ����|���Gz���U+��M�=��4}��3hlL��f`�<p�����뀦��qgMPkր�KTyL�$0����n�lo�ciq�q(=0�ji�^�j&�War���z�3�/q�Ba�y�,I0���t����a��-�pZ�i��܈�*��{�Z�<R�p>��	���ڿ�s���!��V��o'� ����0T������r�������!ؙ�a�6̱&\P�%�l�M璇.���)�/{z��a�X������KC�)3X�
Z�'=A�D݇]�P�Sw��䞃y�vE�Ӛ�;{@�nJ1��)��!{��5gt�1�hdGH�Ջ��d]u�u�͉�!'��abl�� �1�ރ0QFL��1�+)�6E~l�*�Z3H�'wѨ�ꪉ�u�)+
Rk��Q��M���f�(�O�I۰~'֑i;�`�.���H��	�t�bA�������Í<���zy�mcE|X�E$ՙ�.�2���h:�]�HA+��"�Q�N�Z�P��U�;<q4�?^Z+o�{l2Pf��%�<�,U�)j����=�^�ѐսe7.���� k�v��'P1��M+q�Z�8���/=D����>�0�=��}�v����:%��Q�g�H���׷�qtZ>�3Qq�&Eh�a�� �@ �IE5�5�EB������ƽ�[
����k/w�o/�~�W���?J� ��T�'e��M��:�B����q�e��*�>� ;�;aex踣�_-w"����$$<���2�,P����-� �n����b�x�2�/�٣<��GU�<%U`��|�[�,����ī�<,W�H����2F���S�Xw�:G8��Ń�$,�l�L�R"�P5r[c.�0Qp�5�[/��F����pK�c�0��-p����T��&|�O`��Cv7�nw6OB�5�WR�eZ��=�z/���p2��"���v�˩��Kn)XJ����H<��Z�e��½�H���qis2���E��v0 �ub�gBl���Km�N�Z:e�A���vu{����Gwںt���&��^*�K��B5d,$*q/��*g�>��Flo�������5�Z�k@"9 \^��Uz�P�_��?�?D�
��6'X3�VX�&UKG�h�H~4�E4��6�.�;Ȣ��v�z�C�6�z�Jv�Nl�W���]}`���x@����RѨ�c�u�yxq���iJ�V�I�N�_�:hCf���� fb��X���)^����l��C>윾��0[	wߓ3E�N�t�s�U�&(`���|���J�Z}b��4��>���	��h72ۅɂ�����u�� r�*b�hztȐY'��������I����Zc�ۃ��� I��X,^0(s����T%��X��N`U�C]����h�\������[x(#�sD�aذ[R�
U���kuj���y/�}N�KW�Pz�|?��[��&��.2�������[_��k����r8 X$����wzȶIH�$1��f�G{��UM��*�.g��ٳ�Lu"�u����0К1~����W���Aт�d�0���qL���StE�ĺӾ��Snd,#p~����%,�
ݠ���x�_�X��G�'�>���ܳ�Mb?�zm��v�`;��p�0������P󕸽�lO} �4��o�T��aV|�#�}Í�£7r�hU��<J��:�^�1j�ssu�2�
(�6E4K@�$�b�К���m�mЩ�'�Ȫ�I4���j=�v��Ha�;B��<��������>�W,�����r����b�7���٦���R��tm|�J�O(n��_�Al�Z��^_=!��ٸ��p��@!����"'��6!�ֱ�K��-x��z�Y8��WX�i�-� e{�yb���n�禮���L���F��p\�겾R:�4��i��b�D㿳k'Ee�:�M~i#��ζ;�Pq��~2R��.�$�P��cIS�*'�Ֆ���s����:��gJat�;�o�i���2�	��|��dZaR�A��9{�Ct+�^�$ߘx��pl\���v� ���V��?�h�*�d�/&��&t��4ߊd)EHSy��Y"7>F宜����%rˈ�$���t/n�mǁ�%Ё t��&��!i�G�O�����7�����Y����3i?k���!�.HmE�o�<�n�WQ7#h�<�o��P�)��-��nYS��6hʏG|�2\���*g���#`'����{Cȴ ���5�����g|��9�� ��	~�`rR0s���㋋����H���>	t2U�r	
�CHB���e�Q�PXv�>�p}�+�D�ڣ�����_~�*��3�{�X�x��A���t���?| �@ٸy�_�3k�Q�zX��T����`�>4������G����~�Pb-�wD5S?�G?���#�׿������r��e��sn�߇�~�cO�2
/�y4wX�&:��*�'����I_��H�:�E�#4�~:��BDU�9t�� À�'d::) }�&y݆ڏz�L	��H�+���;��Hn��"w�&Ah��%���-���
�Ã�1ર�{��GEi��X��Y�>5\��Vc���g� �A~��<xq����>�w,UrI2Q�U��lVF3�יaj�B�D��ݬ�O]_�&V�����m���VX`��������oמ�;J�s�8�����E�$����w��Y�1Ei#ts�b��:��P��۽�B��u���k�,�z�;Uj�xUx��4b��z�����B���W#�G��y��-cTLZ��:[ҴX�z� ��|��>�74��3`r����o�9�j��f�9�lޟ��uL���]B�צd�=!c~�*��?�둾0I�,��G���8o�*"�F�ҳ�Bb�e���� �t�Zmo�ٔ ��	�V����d�����5�>j�$��Q��1�~���
x����G���it=���D>7R��lQs�(\o>����r�gʘ��ھ�lUk!���m��R��;8�_s��ڌi�n1��4��ر	��;��N÷������d������/�j��}N[��&#�eH�g��)ok�L�~%%�DOa� �F(�Py�[�J,�\r4op�HQ7��?�֨���-���K������QY��t�Z�'���+�`Ė�Mӫ��U����E^����[��Sr;kB�� `�t:-j��F�.HJW�<ه��:�����"�oԌy��~��B�2�	鮁�SG��֎���
x᰻���>�Ch���[e�B�3�]C�IHd=�]�|�i^�����$�5$8�^����y�\��R��s^ژ^m�.e�+�$�ˌF7C�p���gh��_�4�|�5q'��p6���n8���r{Y��I���P��A�9�_���)��6w�����NwĜ���w��8[�n�GҜ�Dm/o*��s>{�\��~�s:���i�Dc8��ʵ������S��H�LI��b�u�al-�T�G�j��Y�_�_�t��s����y2Q
�)C�	�!`u"�N ��4>!�t9ɮ~l�[
� z��(�ذl��c��Wӻ��f�A�p'7ۅ������<��A�.�SŐ�S�)i��ƹ�v%wh�j�,A����z�l9�I|�g� ��|x#�ص��a�X)��hF&LFȃys��Wn?��E��X̧�U͊��H"KЧ5�x��_�ޅ����:�Q��[i��y��q�Ԯ�k��0������^h�xJ� So��w��!<��6��Fj�Q�ěWJ}@�纥t��,���@�W_����gh#�z�Cxώ�����
�r�DSų dδ� /��1�K[��J0�Ћ.:�̓���32u:�xv�釺�ծ�Lt2�����#��M.{�щ�#��]�tӐ	�q�vΘ~�7t\��H%��Ó<�g�Мt�x�>E�O5P����/�/��;z���]�[�L��<��u��]D��+�q��pçh߹J�v-\�  ��pX�pf,�䌿t.�����A��R�X�Wk-i���a|��Z#B�F�2�L�~�"\
ӻ\�F��Ǚ���s|����__��jf��$�niJA�X}3�_A���Y�֣{*0�?���@�kT�]×����ͧ"4�n�k�F�g���'�٭s`ul�M�v˓�r�If��e|Bύ�p�Mn�i/Cn��� ���"�>ɚqq1����2��J
oㄼ<�CӧA^h��B�C���ʏ���d�|#ɾ�������9�!�F�+o��Uc�Tz?5P��)2`��#b�`|��9ϣ��޿>}��x镥c����rn�"�>݈
y�>�p̅t����AB�sDQ�o����	s�m:?d�*=�m���*�sx,��R?��8�.�2�����W�I�]�a��߫/obHz��D��D.\m�lN
~�X7�[�;��*��c�K���풧���F�0X&V����g3�Z�"?��L�/��&z۝d"���q�	џذ����2����	x�`��m։�$����&��fv�H��t��}5/h��5;x걼b�*�0�j�� ���)t��z71jƝ;=���{.k�z+y"摻�woG	�ͯ�R�M��g�j*�?F��`��5L�8E�'��>� !�6��ڻyB �n>S�X����-*���DB�O���h��"4ƹ�`f�VxeTۡ�i�\�GW-�<����>m�xw!�6�(��3��o�?�(ދ�E�ara�RC '��7���b���.��a���p
2�2��)aq����&������CJ���Z� �����xz����[��G�p�{�����y�d�W����:�a�Tqkr��v��W(Mc]��P D� "Tf��W%�f�f{a�dxXh���U5�$9�����{W��Chrno��1O��7y��Õ��e/k�bA�b��G��g��l�д^���:c��*W@�򔧴��]`,��@<s/�ғTχ�ؕ
ũ;��j��\j	ؐ}g��8�5�Z\��?�F�ϒc��X�w�R��Ada3pa�>��qIv���٤0�
O)�y�~���PI�:{�$�Q]i��Tmx�	i���u���0�U���<�yX�9�{�s��
��O�Fta�;Q�V�|�fuF�)r	���˳���Wj�U�B�<Q!���o���)��R����d�뢟[m��?#����V�l7Ϣ��y4U�l���`]�*~M����Z��o�[�ܷ8��9�����Xx����d��\#*~&�����𘟀��w��I��p��Љ���!�7�簰���7�i�aO�z���AwU�_jksй���%&�2�g�g�R�A'�������T��.u19V�Gf��.e��$Г\���L]�2��ӣ��e��p:q�^].F���~b�#�W�ͦМ�?�h��QՆ�V�I0�⡰��kZe��,n�'��=����:M���9�aK5�y {5��� �ˁ�@4����zl���`D+-�T٥��-6F4�!��ߨGnMW�p�'f����31O�.�Dz�𗏸�1�SVH�T��2�6B��Z�D�����!,�<����WAc��V��5�G�w:���Qg�M��rx'���EaM����qe��.���h�d�*K$��P&�G�I�[H�iw�?�|p�����2�Q*��&��4��2�c��-�v�Z�8���2�tI��+�R0�5E]�����%��cK�r(	6e�ɞ�π��)dfjG@���iC�Pxĉ��'�C����T:����8������]P�`C��uJ��=�u�7ԮUQ�d�]�v�PUCF���1���E���s��������q�	����*�e����ޥ~���c���N�u��Ɉl{\���q�)%S�V���t���fсTE�H!.�;�0���qSE�k���9ZV{�7��$�I�1 �����8t���)z�����~�BS�'$�jT�Bt v� \:˒)>ر�I^9��e���t?
!���z�JɌw���_��%����@�K�[��o��TX�4�El��J,^R�!ǩ��Dڙ�S�TQL��R��>W��8U��Y�������?S����sT���μ�Ow�٩{�-�;�º��S݊�F�n����C����P,F�f`�My���P;���Ʀ]�M�vxtbQ��< ����+k8���bN-�o�` 0ܨ��U�F��h��Ӓs���2���d	���T%I��'��LJJ�jY�T�,�w��X��	}����fK�֭�4��,��dԻ� ZX���7j�,R\G�������}q�n X�6�0���r:�"�g�9f)�2������&���az���c���(5R��b�
���u;���h�s�v��P���}�B����u�w�������P�e��I�<���a�����@��IuY�_��2���c�=���,�������l�EN)� �%|�.�q�|�㏞'ʩ�3�h�:����$�/8�Y�
 ��[S� h�%�~j6G���%�� k��ȏ�P��������U�W��AHh��9�C�����9,��n#c��sӍ��{q�uv�;𸵧��M�	�.S�-3�vj�� s�.��P���t��N��1���e@X�R�w�Ƶ�wٞ%V�����+�v
�,�ו�N�,�i*p_`�	X��|�m�It�&��7�O���[B���5@kb3aX�j��l��z��C�q�si�sP(J���&X1>�Rް�:w����6� �-x	L�� K��� ? G3�3�`���%2��8�x��_�Ԯ��wˆF�� � ��@&Z 1�R-+h��%����끄I�T�Dw?���²��{pX�$�k	�E��;^������k? �����HK%R0L�P�}Y��\/�h"_��C��C7v����K6�U#���hSc�r�SЅ��*�1M���`����ܻ�x�*��l���!���f��C��N�($��Y��6߃� {:�N�����kN{#P@@�����*���G�X^3k�a��d��:�G���z3@���d�Ө���R�ܽ�Bt�/���;�ot�{�9��T�|�ܦG��2x�ZBgN��>�a��m2��U�Nf��w�O�|O�y�~��=�ꦞY���^�������=��ld�j���SA7͛I���#�>(7������,2���wI��r����x�}�8��wb�_��s�)k2'��� �M���amJ�5/:!:˟���"Y(�7��B�-$�	Z�����f�� F��Q�8���ڗ����]e�|�ܶ)m���:������⚱=Ĕ}�G1v�y���[�M��2��|)����P҅��b ����4�br��{ϳ7��=�]m�x%`F~�?�扃y�}�^V����5�\���,���g�P��#�G��8Q3�S��{Q&d]��XD�y?<��!���X�X���o��ɹ;*�J�,�Z�}�V"1��5�-��U�`"�5�,�kS�rxuvM��f���;%yL��jxE��1y� SO;m9�w��h@v}:��1]?]M��⹂���⃉�T�n�U�ˎڠ @p^������H�ΰ�)���(�if6��#hr��U��W�U�r���U�I�pK9y�0��0�ƃ�i��{��8��~����.}����T
�c��-�z���������H`COG�&�y }�%���K<w�d�!�+�Id-9�X�X8%���5ň���t/�O|c�<js�{q�a�
W���[� ��vZ0� ��}S�\�.�Hg��eL�8*�]wK{ڗUeo�1M4�0w�Ti�̿k�Ce9m�s�;J�X��ٮ���0�ɱϲ��\�A��gWˌ�Ã��/�eP�������Tږ�����P���p����Ma�B�/�/��� v�#��jA��X��-�L}�X�3�g�8����D܌@{ZȗV�U��?�9�=u<3Y��8�Zp>��[��r��RZ
�����F�[��o��g%
��/�P :��A<���"'��A�����0N:�n�v>Ő�^� j$)�Tgb�W�Z�?���Qg0�r��}M�w?��@Y�3R��'6V,�B#���7L�Rv��.��8H��+����f�8ă�a�3/���2�~�U����c]�
�w���CL�t�w�-WO%C�����_�G���`�ՠ�Î���@�23f5���S�=O�"�mh�Ks���L�q~�$���|�{ U( v��?Е�UlX�]���Yq��r��i���g�v��v��w䃓(Я ���^�o�[��g����z%N�A5��숾/��k�.ٲh��[Ik�i���ko>	��ݽ�0̎�j3��Q8̶����;�}$����!F�$]��ݿ�-j�6'�-ҡ+>�rI1*o'S��O[L���_�\1~�����~�.'t@��Z�H;6���Մ�46�:����d�ˆ�<��y��\^/8lx��\aք�xaZ"��ӫ[tlLy��|���j�.�.��"��@��%���Q��,o!S�]H;@=�DP'@#���)��~S�;)���k.L~)�D�^
�~J*��;��&��y\�$>�K;��1��ߙc��cGb��E:��"\�z�KN�12BN�*� Ѝ�V�]&*���jB��h�2���b�?�a�3 )�m��� ��� T��j�������7A��B���x�[�?p����&�RG�՝a��y����q���\�����$��vA^j(��[c|���F��Б���ک�Y�:�l3��V�>�9�;ʵ�f7[��u@�`]���YO��y��s�١x@�<閇�2젉��q���LxǗ�·�hS7c�ײ���:�{,@�b�:1��rm�q�w��'D? �)�̵�s`�߹�������Ee)K�N��7T���3��x��w��Xȹ��8Pf���<o�h"����	�!,}+ݎ�|�Duק ��X��Y�K�/G����g��� ��Fח���9�]ae=�o�x!��]��$�Tzʰ��P"�c����)%5��S^Y�Lp���@��ܐ�π��"�U�8m�!k3�����Y�P,[���5����3��C/�˂c9��ē��a���y�ͻgj�0�T�4�`)���OAY�Jxnb�,6:Ήo�K�r��C�����%�p_?S�Is���m�P�����=1�b6�|��נ�u:����*y\6:�,�4�^I:�ë ���fV�߼���Q�Q�u���b���xAwr��o#{,C+%2�d׽�x�ʰ��lT�
(4��⒃����;Q��4��G��C��L����.]�������i��ѾAh	�P�f��\-�>�o[����ug��\?���Dɋ��p5c5=m=5���L�Ҷ���s[1;�s`%����pm�����> �6�]�d��~1�)���uy�������������M���t��e_:B"��:&����>Jy̔��91d�G������	��+��.��,���s�Dy�n�d3y�QNK>��67 p��Ǔ�X�b���l]�9Z�Q���;́=����
u�[�pJ$��@&+R�3�	v�Br�kɒ�q�³Ik��C%4l;�`�����Ur��v��9��<��M��ذ�Im��Z��"mcE������Ir�������`YNT���k��萦U�=�j����������C�w|a~Sc���YIE6M�0q��&�Np���\����N�B��`;�����w��˧=e]g��L�c��N�B^�Ӕ��@����`�Rm��]���� ڤ� �c�F���w������Ã�U�si��U6]�}f�\�� �*{C���5˱�K0��Zr!�p�{n<E^�]��5;��7#�:��Z�]���g��ˮs>Y�*r��L�\�f'�C�Ƈr'�8�
 ���/��K.�ͣ�	lUKzn�=,]j�M>�a1{�z=
�91U�K���itC���%����S�fίr� �)�'z�8e�Ohpi��0�k`��b�6p�oO�)���!f"��"�qJ�d����\s}��"�#IN�k�h���\뻲�����t���	n�M˧L �� ���ݰL_܃-�#�j��.9�QL�,��Y恑;�y�m��9Dn���gx#�S��0�]0nٚ��A���G�:a �>� 9I����M���}l�I�p�$�f�d�B��2I[DA��?i��c����2@A3Z^ �m�>#�G7�&�a�9�Ǵ�M"�׸h�[3]�ǜH���IS��Yr����S�f0������Ջw��X`���Kr)7g��_��Y ���=�	��8ќ@'�:���bn:ED�������v�+7���< ӯml�E�aE����*5�-��ʳ��/�\0ߗ������A��ugC�qp��]����w!�/�|�(�U�Ń�8�<���@�r�o��>%����}��)W�/UD�?���k.n�fc���ؘ�ǥ��ʹY"p�ey��q?D�L���y�#-�k6�v��u���zY��������W/�$C��AA܂:���b�w`�L�7�%1/z�Y�|�-2�]A�0�n1O�@N�~j�^���&V��x��)�=h��&�q��Y`� i��@ͫ;��٨(��t��j2 ��^�{��'����ն�Ew�`6[r�Ŵ�+� �9��5\.><.���-��w�0q��⶜V|#��i�K��ee(�o��]Ԟ-+��{fdV��
���e�� ������֛xR쒫��!�t�f:$x_ᳪ=�c�g�!Ш5����~7ٳa���-YQA�|���Ӄ �#��
��=�/��k�C��ʀ` veҵ%�Hq#��+�5�8L�3�������I�: M�3+Q���E�6]�p��0/�$���mؙ�9���]K&�j������oz\���Ɉh���	A�I��φ�A�4hY��.Y�X�U���yF�M�;kFώ�]����� ����"�����j+�c�]�M�I��)t� ��b,�v��0&��ll��L�%+�b�	��ǉ���\ю�H��[z�B��-�Md�_mj�٨�h?9[s�b�%"�r����s�_wЦsrxN�C癤[})֓1j�D���w��BCyc����/��M犩��M�O��!p�ٚ��b�Ȫ�dIc������7II�1$UBRk�I��#���ڿ��yH���O������v#b����>W��'��i��M��c~�uI�j�T�'��z�;1����_0�T0��+zX�S�� �������y�`@;_�S�%#0P��_�R'�P��wn�(g}}��W(%[b�jFL�ZcQ��,��pP5A@u�b��&�� ���;��,M�׬�?��g֞��Y�o��0���ܘ".��O8�xi;4ԝU�(1k�_�Z�;�{݄�'&B�����eq��c�h�6�u'e�}@3Q�b��h�,ԛ�*X���.�.�NmE�K/�.�l���ո�m��V3��������f9���C���w{{L�\.y�W�}�ͷ��}|��)?�D�V�F���dP�*�:��_�Jb���7�7>'��Z�u�ml�O��u^x����F��m{�=c��`?���?di}=�Bן�7Y{a�`�%ic@���K�=�Tf$![»�3�d��~�e�_��x��H��tB3�&W��\�y��[��������f�@�ƄHj���0KE2kF��~�~+�����[Zl;�zk�#�n�ߗ��3I�A̬��jc�-�Z��I���m����LX7��g�A	M�*E��'�~B|�����T��!�?L��� 7K�S��݇}	��s���g#wO֋)�#����]�� 8����f�s�溉�vsf�BC���1�����B��]J�]��i��)�
U����QV�%����8П���n�r���	}3�a}Ll�]:��%+�K���^��|�a*�a�=k3��;�@�B�Dw�0����*e��-�bS�v���ߕo�O��-�k�-�]s,�g�j�Dަ7�� ��Ƚa�u^�w�h��X�jE�!E��������]0'�(�@0�K�׷x6� ;g�Ψï]���c�0���Ȗ�j�����Ⱥ��G�I���J3AD ?YE�ȲF�n�xrd�_6{:�����y����=L�c�A�m�kQ��������ϸW�oF�����Pv�f��{>���*Tu��N�l�GȔoGv����iM���9y@�����=�W\�(m���]���dُE��j{�M!� 	mAv{�G���ot�F82�����9t��Ո
�@�'�ϳ�X�>G
LA��,E9�ʆ��gi��DHC~��Hp�q�©�pU�?f�!G�?����q�������s�;*�L?7^�=�BMo��aC)�h*NHhǫ�HY��f/�g���)B�dh��FCQ��姓+���{xg��h}��i8��P��\`ǙF~�[���E�^T���j3v�r�ZdTX&���%��Z��&��W�~�޽N35_؎<�e���o�¦����PT�<៘�xo�"t��˂;����1#�܀��Z�cs��`s����k��O�V����k+J� ����
�Ȍ�k8H ������b%��+�g@1�#�}��̭�� ��*R�{{�o��SI��]$��~�bT[�cl^�X���ڏ�*���2�Ϣ������!�q��Br�/6�?u}�`'���<혉]���X�:�m��'kx���6��cE��r29��z����k�G���Į4��WT�|]!~����'�.�b�d�\\���<���C�f>�SzQBp�F�j>5Oz޷P�b��<��4�`�8!	FK�9] �	�*r�����I�y��kߒc�=?O.�|A��2����s�i��,��qD;V��ǲ��P�b��؄�p�w�6��Um�j��D��I���\8dӂ�|VE�u	������u����$�4v������Ʃ1J�} rH/ӛ7k]K�ȷ)苜�Gm�����G��u��˵꬐RdV�, �^�jE����}x�Os�Nœ�t�ab�޿�#�"#&���7� �GA��zi(�^�<��;�U��0������g�rp��c1ed=��-:��`�S��: 0�F+�Lv�ş����<n��x쉑:�����~�Yd�]������Mr ��H�/_���58����<���-��u�q����y�	B8������r���ZX�+ q/}���O�C�:���r�,���o��˂h�4扻�9��bݢ������1�� 9��A�� �A}�ʘ5�ڜm���$@+[J2qp'�����lRV�*��t�o^��OO�0��8p[jk)����5Mv:_s�L�CRzD~����/��i�7Fu,x;!CO_r�����P"->�HCla�AQ'�	�7�a��=�j=9L�(�o�F���gX�'d��;����mT����Fg��F�'��rBA!o���2$b�V��Ez��<d�K�"5%c&1m��Ϳr�����a?��#��u��Z��P���F[kz�_�3�[_��9�s��H� �J�^>oN*-!�m�cL�os'��Z����k��(���b����Ҥ�[#y7�����8�G;r�T�9�!k��k��&���h��eB�4JH4���utk	h�_���gx�nm�4��*IE��o/2v�#���ʭÌ�Wya����c�q�f �Go���kI��UQpw�7�a����pd�w��>�!�Gӎe*a�#���EeTY"a��'O��v@?�ګ��eޏB�y7	�E�	���l�1ϑO'��2��s;{p����i�3�'ֶ�:�}5�l9&@hgm��i�{t/�t��x�i[?Ct�����X,WlEY��+��k#��Ynk��(=�$�7Vkj:j���Bc����x��W��v�����8�o�;�^�v��I�б:�f��!D��>)e��V��3��/2w��}�B\33o�t�.H3�Y<Qߛd��y�e�|��m����%l�	W$��3�.{�/ [k��cĥk�a:k��	�@�
P�GД�a��ϸq�8�R!-<2w0�*�p牁����S�) �	���BL1� �vD�9�Wh��Lw�+B�qaO	?�IM)7a��*j����('�!1��o�!��Z�0�L���;���Q� �k�D��{z�3�#����4�C�G���hJ����<ÉxS��#���~_��Hbdc�8������y�<�b�V�9�ܕm�TW�i����aw	E����t?�<�L��7Q26G��L��a]���EH�����F3����g����.��3}��a�x�<N�AQ���м}���N���L�*<*\�x����x��p�7�5��:۲a
�7[J��HP������,���Egx�[F��_�H��e%�e�)r4�����aU�#C��MA�����]�$2�e�=�>6�̋;��5Q]��M�	�`�oqP�Kl�afUB�%O=w�����%)�v��A��D�3�Ir�Y��	�5��!�G%���f���H�N�l��B�H��t�ǂ�+��Sp 0��i|�7�2M�U�NFn���7�n�?�`�B	��������QYe==`�Wv��O)��܊��h�`��sF��ϵ�$�_�nW�Ȣ��� ���Σ�'?65�|������I���*���R]���v ��do��t֮�ה��G��e�9;1pm̩���k�W={�ń�UJN�gs1L`̼C�׭;lղ�/Hy��D`j"e��1i��($6?@\L�h�v���Tu��o)�z6{�^K^V��5�W�2�������y/�2ԇ�C���g��|5o����U(m�ܠR�NC�WC3D[)R�(c�iS��7䫎7���E�(�/�:9���ŀ����Y�dSx`����	�~�9�����AR�� �JMfQ5�Q}Kr8�}���!�_!<����9�?��XU`��Z�Hd,�?�R~i�,�[5+ٓ1W9��iaF�D�}:`z굶�0IDc����z���}{
i�S����
�P��Wùx�ܛD����΅Ug�fǊ���+��~b��� �̲�T�jR1f����j<#/ӛ��	ȭ7s��hwߣZ���k���eV�@�����ϔ��o�BgdSMC��s3�TF��C��OBA׍�NG���D���O�X��R�����dq�-!(�p�E�|�"�<FYv�B#�Z���G��%�!��~-��nͅQP��a�FŞ�V�yX��V�
���{�A���Vi��A�zS��^��w���<*�\I]���Ƕ�5�6%a'�D��D�#7f�YM=�f��ROY�Zu�dI���A���\x������@
\	��z!陾RaSM����H��aP1H���R�:,~[��2�g�^"!���<^���M����(���i�Uds|�J�<��U7ʳgH�M�q� ���6Y"��!�1M�`�f��Q�{��>`����Ioܿ��>��UB�>��L��f�[���E�\6����#�,������k�H���a���!�^�ɜ �= ҝ��1�_5Ooi$Qn�9�	�IeRXZQ��3�?�Fyk��/
j -~���U�Ʀ��3l��.�;E��:ݢ:T��h̓w^�[ܶ�7H��w�.���4�<U���znn:�����2"�{F�P�£��-�H��]��n���/ؖ�?�J�eg���D�ί�`��*�S�ا���y�k��<c/6�#H��#Z������t����9Yw�F1��РGq�D��rK_lT����gN�a$+�2A����U���"E-N�E�>��x�����⫝kI~f����&���GG
W^�r6j���)V �Ԭ�D����~�08��(�ˎ�ǁ[�m�ے�f�02ޝã��p��c���"���y5��_�đ�[�U���Q�0.�}����'� ��7�����*��N3���������+�����D� G�ǧq	^�f��~��<k��A�X*����&T��۝-i�-j2|=l�1k��F*"\��x6)n}���?N!��7^�z��9�ԯ��NN-���xK=*qBy�%#�<��X~����ٟ|��n��x����;����?pf���j��/�K�|{b�Z���8�pn��l�����tz�XG��XX�`���[��p�,۶N�k� �xؾc.�g����	��:w�uLؾ
d�V%L�M���Y/�W����)��_K���	E��3B	��C�(���f�ޔ�:������"��~Kh�,�x�@�������G+q�t;��Y�-4ݙ�Ϥ���	�{,6�@L9�#��m��dFT�/U}���:�g�f�L��x��������[�2��J����H �g=�聮��j�w�� N ��G��aG	hq��
,�_s�s)����(Ȭ�W#�~3���WEk*�]F��É	�6)�vኟp~֞[�	���P9��S����VQ��[��e�k������KYP�q{n��a����	��<���ԣ���iKꆭ����9ܸ\�4��@�1-���5A��4� X�/$� U$K���{��Rʁȝ�wa���P��� �>���=)f�է����_�-�����[�L�8�נ��s"�h�"�D�~+��`7N�(�F����Je|5q.}�E69 C�]�mL����q�z���a/�	����4&|w�K�Ob\�̅�+����߂���I{Q���Xf� �H�K��/���6U�;��@��+W!./�+Z�%�k/�6����M�Ö��H�M���㯄�b��*dJ�By�������_�����N��ٮ��<2�n�I�@�Po���48�"I܃�t>d�os^�Z��>�����s�b)��v��LK2��0����L,'�wo'���7�K����A�9%�8Ql2��16�8��Rc��)�cSw]��8s��%�Xt���Lrֻ��>~25�u�gp���Tm|n�7a�ů�\���&}�x*�!�F���4h>h�Xp
	�����+�#J��c��|`(��īⓔ�f�^�@dɼ�ؕ	͞ϳTx������ ��zil�����q�t�|$t�4�l��]����7�r�v�ED8��C��2�^�u���za�uL��E�w�U3bp���3Hk�:L�.�	�M�)���f����Ď�9�����q�~2����� m���!|��/�J�e�n��+�(����		�኏���c�73�LA���hgI%��>h0�wлH�bq򁱔�5�����LT��܅V+#	��B]�*�L�Ἱ��NϠ�;� ܔQ-�K\@���?pN�.���dԫI�M��@"713��Nr�E�{��/��	��۽*�Bp��{�b�.��q�s8��:��[5��@���Y\�������xu����20����>m�<��?e�!��^y��>�6�x6?��K�gV\�+N���v�=�G'�^'���.��}�W�АV}멑�g���M���͔��`ǈ���,�b~]�~a;�p�hia��9�=�=�u����t�̎�����#:���� 7�2�7`�B�J�n�B"iM�E����S�([��!^�j!�4k4������K�|��r�S�����A�9�P�ґ)ט���u9����*��c�hC�d���I_���
ɐc�̕��;ƅ��`�X����M�#� o-=~Dts��z�����%cq	��{rDO;wĢg}a��q���/ة�h# ba$�M'��&����G^Zj��8y D������Q3�d
k���tQ��&�(�$�'��V�^ƹT���:�*U��r��/�Y��w��	�}+p�c�zo~�y��[n�c˫;�6�-�^<���s��ϯ`��,�=vy��7�m�˅2��3�>�̽A�ܩ!8���0sF��Ǟ�3'���L��;6 =��"i�L9"7`i�A-�}�۷�1�[ �����/�/�#�ijW�֙��Q���s���#po��ݩ�oRύ!;��Տb(Z3��4
�"%.Ʒ���T��G�X����p%ٵ*&"�*
0����5��{T��5iIȒ���6�������Q!�{���͝�x)KJ����+�v{��7�ey��I�Ҏ{���ͺ4i����f�_�d�.����Dh8*РPѹ���G�����>��޳��_�3�G���o��<�;����k���dI�>35+�>�M�XS����] x%}�AT�<��g���8��2�4�ڪ��dc�ŌM�$�����M7����3U��
0.~- i�5<�zZ �B������[r�RF�8�
<���T�F����p�c8�]~�+��'雪���EB @3��S6���S�9��me�v�	��r�� ����1�53s(Ɵ�M��g��FR �I;ւ�(��Z_��s�o��=�O��2]�Na�Z����!a�W�)<�3�=$^�5}�&9/A0�˘�?HM��Mͭm�ڬ��]�'��@"n�rv��哙n~f3�B��y��m��҄4 B���4�D	g�*�} K	Mu�-�BQȚ��W�18�xP��Cvx��61���0�yբ6NYbBN���&����@k����o�j��������},|z���1��b����e=��e��k�����t#������rC�ߑ�%>ٚ�;$�+�Fo��L�(��?,�XU�"V�`[ ��>U!,�4��	��N��������*���'�w��%Չ��Z���{s#o�C�b�mA��d�74�֡:By�\��
`�����矈��Õ�^ z�aım��r_-P5���e�y��/UE� )�A�4�"�}�<]�P[p`?����o����߶�0""�&<�*>��9���y]�k+��[��F�M��d�,t��} �|�(����דZ� ��I&� I��U����e��?��B�3�;���8Jh��]�0�ӭ+Ė�G#�@�t@4���̈́��B��E�v��k3�U��k.��WE_�G1���gy	:�Xc��{��V;m�������gd�y��E���o��-y^��U�B��t5�w�cI���IS�\F�b��r��Al��!#�~���v=��-~��M�?S���)lj�k𴧕�}mה+��>X��8ܙ?�.��_�%y8�	#�I6�x����G�>�����S���W��g�*W�[��E5���S���c�54O�!��K�d?�;�ɖ�(�Y���P�;L��uc��������b5^���a���لcB ����"���|�FrH�`�����_�����5N�Q�)���*
��Z��Y֣dm�*f�>��x��@�+���g�ukX�r}q���������l��6���a˯&�Es��xw|�� �y�v-���0�ޡQ�UL���^�a����t=��}�g��V���|!A$�Q�<�R�|��C!y�"��R���hW1X�~F�	T(GdL8[�e�:�U(%��2(��]�ֱJ�Ss�(��t�j�0�� ����hcT;xͷC틍���� ���Y25i7v�w�K�>"gI*�W{��Rqΰܴ�����ύ���Qǁ^� �?f�"�t>�CWۘ���`�N��D��됀������[X�������(u�)��w�>�������?�TE6��>�^����cSᛝ7��3�����w�,�Gzؽ�k�P�)���E��A
-e�����͋���R*�sf��i"�l������;u�/���E��)��[��5�s$�}Z��'�8������h8q-����7��	W)��$qu;�V �l�ϊ�
h6~���#P���.��օ:�X���� �Ҟ�X�q�����n��\ KX1��k:�٬c^�f�b��A=�.v(��N��2��9i��D"p9ޡc��2�@	����eyZ�ވ�5�M:�$y�8k�ub�vG��g���8C�'k��4' 4��@p`�c=˩�E�01�A�rQ�֞c��d�@��� K�Ň�5�~t��%���C�s.�t�e�"J�[e����KTx���`��g�D�J���D�]l�D���y�]u���r����u���<�H�x�gON*h-}��NG; �WR�4R�}�&
4�c��H�a���(���`Z��Q뮍J����n�G�e��.���sQ�x��h^X����YA�5R�I�h`����8;%d��u�՟R?�e�K�Oq��j�gf��N/;���㭤��$����p1?ė�S���CY�)��U����ܗ��2������e�C�����|f;m"��;�ag��t�z��c���7���Ih�Fl�[Qha�T�
u��}�^�x�n�$����Oad� W���U��l��sg��$P�yհS�8���M��ǹV�N������e�e�Ak?���"L;�,{��S}h+L��(5CPa�k!��#�#n����rJ��������!H��3c���I�T�>��P��V��tMM ���)d2�{��2�+.!�j�����L��I���xc!��U��57b��gT��W���#��ح4A7[I�7T!$�8����[/aK�æ�W&m��2�������*�?2�0�$�'�@)�t�S�(��Ҫ�7k��%��+��GC)�~,ʲ�֢"�3��nk�����U�_(}LEy�I:���y��5]�C��['��z����G��dG�B���2K��6Jj�&]}� XU\ GN�����k*�n->3ZM��]%�Qw�h�>�n0Q6��y`	��V�F��p�?���_�1��9j(��>��S�G��)��G ��q�3B����v����r�ؖ�w���- z����➁������\��6fwZ#��İ���|���N��^=�SS�����d�!���E�Ӟ	I�$�0�z���ۚ"�<��p�;�ņ{&D"��Cw���yatƧBnz�a�S��vl���Q��U���4�@�-�(���-�Ti�H�����j�{� ,Lᚰ�Z�nD����L�=�ŔYcOT"�-TJz�<t�+�u�3����9��)2�R���̈�(�|;�ܪ(_Lzy���h�T$N��~P]��d�n��Y�����(6�O�
'��v�w�GS�X���T'��A��%�ى��Ob�6���fE�4���rUkƉl��KQ�܁�X�"m_K�{�Փ�O�����e`���{.WŻ���E/6;P��[.wL���LW��H4Ug惷����/�G�1��3:�����,����(�>=��Υ^��ұq(�l�-D���H0��"&�,��r"�(��.���ɡ�ƹN��Gc֖�=�/�Vho��t��.ێԑxxቇ����ku�kѸ9���u3W�~�?��\0p�E��3��9�P������$o�<S}�0{ ��T�a�i�O,�F��r��=WLb���2:��f4	�D���B~�^��s���U����A(-�rq��ٷg�K�w�t�iQ�4L���G���1W�%eq_�W괻�~� G��\d�\Jʖ[N	# ���8��H��}H�L��S�0�Uu*�YD��%�f�+b��a���+��A�k��l.Bk��7��������j�a|�AƲ���;c��ô7��zb�
�U|d9��Ȫ:/�h��g�g��Vt�W��"�t��'"�:nC/\,C�t�߅<���&ȯ�zs�<�Sy�\`��L�4��	�C	�f�G�^���/5����'ݔgc�@�"��}��7i��0H,CD�DW�p�<����[b�{���l�N���OK�� ���i�A�^��rޤd��avqu8�JRw~��Q`�~x��u��h��l>j�ғA��(�6��]�iũt5�q�ή������Z�E��� Ƈ>���~��qےZ�n��I*�u53�p2�3�Gv��(4RA����&�� ���4U��2 I[Z�:�ᷦ��@D@��PVr��Ȕ��FG{�6����^���
'[����+2�W��n�#~���[����n/�ǲ�U��t�1�Й���6KB��:Q��c���?�*	o���g1��=������X�O�y�c8��Kz�h�q��<ǅ�^���퇎��\�[d�����3C^Qn	�:��;���{�3 -T�����y�b$����"�:rs�#����C*ձ�����q.4S|�F����K�����~T���i�"%8��
�W��F�H*�9�]�! T��Z(���n�ڪ�'�wta���xk'������&��A�f��;�.�!���KG��2�F�6��;,t�K����*�!��Goӏ5�?S�-�@�����z���	����*���j���}�醳膽7����(j^�V�#C6S��ٌ�� ���������|�l��b��vC��s�~��c=
��M��H����mߘ�A��,��w>�U0e���&�c�[Y���@w�(Ę�t�0�joJew��'[ܱ���z����IQ	��$����kTt������DaJ����e�4�$����W�A������5�o�� ����F�_S/ޕ�򵉠|W�:g`/ۏ�u�Xu�T���b��ﮈ�P��7�����_&���ٵ��dߧ�}����(0�US�Y��v	��as�_8ѱ�-���̈2y��`����5��[�`(���kW����>���=R�����y�GA똒O�Ǐ��]`,*�-���;�A��1N:9��Fݝ�L9��nrdUG��w��=� G�\^���j���>���{�l���
����xg�~�w�P�D���֞޷c�2��P�]���oD������2�3tY�>��@�=��f����������xj�L-D�����C�I�8&��;�&�q�WE���Z�Ģ��K N�u �����X=J��n��1;��s�b	�
Z�� �����-�� ��[�n.�ڄb����WIhJ*��;�F���N�xҏ?���6޲'�X@����l�+l��ߘ��	�G�p�_����N��/w;�6'_����<XJ��	��x�Ys ��ƍ�,�
/9��=�pY�#IW�m�=r\�׹���m���[u8��������My"v��i��|��hna �y`<r��Ps��ĊQ�҆��x���������X���b
�mu�ۭt]]Y���-�h�5��������z|C��#kԋ��9���d��m"8Wd`hz��Z�u���x�@ �o�H\H�yUU'�U��sg\���S��z����g H���B�c�po!�_-V�? !�(P~����g:�E]F�Q������T�1��
:��'F��� c �P�\���&W0�U��.�z�ݔ+�}:�^�~>Y��I����}��{�}�;f,$�`�hY�=t���n|"���t]��]�Ԏ�>��V��9jx��{��+D���@,�e�P�_*Љg��wo=z���/$0�ئ"�]�Q�WߟRoOxg��8P;��:|�	��C�& R�\%�O��,>&���Nױ�rQCH�.P�9k'60~���g+nV��!P��e�����X�1�ٚ�8_�j1��c7�'�e;\� g�$�Z�b>Xo����)e�윋Ϫ���dΖ�a��1�%C	-��Փ���4װ�(���8�#� FS������,�uui�^��t���5-;�Wh���@*�������&b�ǵ���i}��.�W�a��l���xB�|u��zI��\�
�,�1��ٗl�'�V�o{������	v��AFwZ�ɾu�������{&L���h
����xF��ߞ�X�5��JW�E�kv�\-�ڡ�*�Q���a������lR�L�E*�׍���r�/��N����`��X���A���?�������5l#�� ����a�($����L��x�2���а��^
?�@�P��3 ��>g�zM�L���!~���|	*tR�`���'�^*��wm�|��\��$Zg���b)�s៎�
o�,[I��d��s��gP����nQ@?;J���Vi���md!��EZvŮ��u�Mj��07u���P���{:£ˌ����l{�kj�e�Ҡ���$L2z973e�C4jw�k$�q�6{醙_���v����p1�;����D�=T�k�"u��GUKT��m��Kք6��п� +�s��\/�9��a/D�L�`w�b�,��%IU<��@�<0��r�C�Q�S{?5/���y����!�]Εrom^Il���sP� /������@�V`K��mu��I��	�^�̅��AX&�n�u�ww�M�t��� �5��J>�g��^�W)���3��{	lV>݋T��S%�s�/ 	D��L�`�F9<�wjl�dk
����2+o�u
�����0�[��n���M^yϸ��M25|a����%���z���^��H��y����e��K(9|��Y�	����کS�C�-��,�?��x�ʝ%F�HO�q��6<u��]��⽽��ͫ��fL" �=�ɘk� �4�>
�NK`j˾��0RV�؞O��	\�3�"���c�XÞ��9���\�Vu��bҢ	2����4���8ֆ����i9��O��ŻZ�,ViG�����ޢɡk6����DӸ�����$�s@������u�

)-������FY�b�i���ǹ���i�Xq�D}�Ԓ�A0�e��d=M�QF27��P�����c�S��|� B��hhߏ��4me6lI2��	w�i��|VP}���iEnx�s1��G~$g� {~���f;2��P��^=��8;�w�&c�=ɨ�����J�%�W���o���D��;���O��B���Mk\.�u%T`��4u�h�6�d2g�xN_(��B����b��Bު�uw |������>��c�_�$%�R@[��QU�zJ�Ky4
���SF��K�c�6��|�w�\H����j�v���߂�@G�.�鵥�����x��*��&+�E�q+D|���-S�Tٜv�:PQ�_63�E�[���N��L�\�N�|��{MK�W�����X�%�?GDQZ��䚒;��?Y�����E�XP��h4����!+uy�H� ��Ɖ�`	���a�n��&�����_W��"�h���<T��$5zH� � bћ�j�yH�]Z�5�����.g�mQ��\8���� t{���ٗK�Xp�}�,���ox]���w)�6��9�u3���q!��j�譫�i����`��}��4��e3$qhCy���pľo7,�W1́��+*�f�t�+�Nz~�J�ЭEP�1l|���gyU�m�w���?�'U(5vW~I�S�%��mt�6n�2JR�6�����X�n3�k!s����f����|'F���q����l��5��Q�K�@�H�I�`�.јg�aj�9X�@a���p/�����%C�z#�,v��W�����܎�Q o��Y�-���[Q�$KO~��0�y�ZVd��_�\4N�1��/
�w����ց�v�@�Нr�@r�S�������705+3UD��M����p��g� �S�H�>�ף)��g����\K����<��[(P�$e��r�aplb6_љ>O��Qv��i4ښ�;��K��)�U�1wc��L(欶�D��>g&��nE8��-��^8T�æ���A�+_/L�PʨR�Ų֌_pSE7�O 	�^o5LfWi�O��R~q��|3w�F���(JՔ`�Ȱb�_�VI���/a]�5 ;ON����DM:���k��sU��C���9��h)��3X��V�����g'G{�����`��I���5���ݦ�:��6n��o`��<�$S��նGA���((ْ+V�������+�|�V�uZ�N��W�n�H�x.�;����������2j&�ڳ��){J�E�:3�Xs��_��kJ�9�>E�]/�X{~�&�D64./~��gE�Ѐ������M@�o��:��(Jѕ�=9n<�<�FZ�W�ר;Y4����=��t�跸sd�	���u�u���}��~$t��N�SD�_��O�'JC��d#`�� %�a�S���3����i���9g��_�ݻ�'� X���D4J�^�n��j�͓�7S��o7��*`�KN�F/㒘�,o�����| b�~)7�ń��7,�C@wg����0Q@�h�����9�\�����ѫv�<�"�B5a�l6�U�r	���D�Q�B@�D�;�g��_�N�}s�K�7lc#��curS�i1�I�?$3y�0�%x�&�W�W��6��ܐ���dmY����t�lfx] m��g�
KL�S�*$اQ�p�c\r�jU����`�.�2�1\�!z����m���Qx�#�4��N�
L�I��9*�ѿ?�V�Dfiٓ"Q�?���n�@r�m
��_�[̬�Ɣ�����T���O��E��8"�x�v''��8�m��Z�̀���Z��Zi��8����y�OD�u�d֧Pb2�`��<V�Y6�f)�#��}��xO�d�P�C��^�W�˥����W��o�٘�e�0�x�����-������0��RSLx�r�=D�Ps1.."�pdi�C<^�>�4%gEM���#�9����K�]����M���m�ؕJ�vJ�����/G$��Pupӊ�(W����<(s��qR�eP}r�6)���ô�j4N�K	~E�p��Ht�RY���-�c�/�2����?7)�3U����\h3�^Ո�n6�4�=�~HS�K�`/�	�$�j�ed�ڽm\j��+a��^4�DA��<5��Z�;4�}Bn~#vZ�u�}�+ ^���ޙ�sA�htݪc�΢hL(��wç�E�@5��Yn+$��UN�nn���j����!T��k�A	$�_ڽW�8-&�
�W)wn���g:Sq��G��1�)�=��Q'���'
��&�_�֊�]�2�M|
q��dn��35� 3�dP�t�>�P�^�Q�)� T�!��5yrz��I�~~{�o.�������홷�����F~Giڥ��8�fKXm�{]��}�O�r��!����HI���7ƖJBe,骜��a��ކ���MS0��Ik�lV��4��k�_� ��n=�d�'-��a���X$�?Ǻ�=�&\jV�p�C{J�?�`�h����p|RK��Bj�d��w�쉰�D�u;t��!�8y����l�56��iMA���YU ��5$a'sw	����׏���̹����ǚ5�p�8��������A$�T�n�F�F>��<�·��rQ���5��v~�TaRme��Ĝ�D�����@��e�K��A�$�Cm��� EN���6��}F�����H,�/�_���{��L�z��~\��Am���z.�^A���횴�|�f�
�4���J|o��{�&h�O�eW����Ee�Զ�ja�*�~��_�D��s>���'�dw�B��U���rEDdU�|0���5X^���0J��ޣ�/-�t<�t��*����/�*��
������vp/�U�ֈ��a�P�w�#�0��y�-�m6��iG�{`��aHH�X+�6p���YIːh�V���`�Y���V��s�+�'�-�ǣ�+�6���gM��r�[�I�V7.�iv[p� �#�����+�r����=��!��ݮ�-�OD���s%�c=��R����M3����$�p&�^���P0d�t2��J'��'|�>��Jn�s8�O�oI���4r���
b��Ȭ��,]�X��^E�� ��]K����x9<�_J�^�l��[�M�w��э�%Q7��������kUC����X�\j�d�*�A�rX�`����)�N
H�J�<|�c1$+����N��̎@δ4�(&�ZXv�*���3�w��N�a�t����v�z�wst���Xn���@s�Z��;~O�v���J<�.�$�Z�`(�ָ,�ws?��ҧfq:qLs�Ae��l�%�~�D�w@�	_+��_Ckw+'(e u'I$6m��p�7�u/m��|�1$�^��v�D���l���\S��Th�"�m����cl�_������a�?����:Y���hL+��.>�=	��y�`�e���<�"��&m]nI��i$����X�!m2v���]I����A�(�q4��ȁCA����#(�/�X�?�K,"K���u��[|Ӱs�����&��d����������S�g�	�H7bO2㖪�4�5���b ����.��g��*f�ۨ�yL8qq�g�����#Z��9T�-� j���2ﶽ+
K9�C���W��xF��e�y��ȢTŪ�aj~�	�=r,Wp�c'�z�����g 	��̶D��I����_X�s9 Z
�I�H}��I�| WPx��ƻ�?m�i��(�&��"�%�j�_\�Zt_�1g,��[��L��ϗL N��4���|d-y�7���v��3]�c��w�+
�x�v��7՘�"��IZ��O����(��Ô�Z�i��(��-vωud����@-5۽i�z�����h�����p1�/�鱃�e��^�� a�&��<�������R�vN��Ό�7��/���J�@���,�Q�r�p�|֌�)�������/�ޤĻ��ϰ��U�ࢶ���6�7rY0[78�l�\��%0����x|��*�[��ٵ^I1�P���:DQ���3�=���ߠW�����������4,��%��n���0MA��|]��	@�h#�`�M��詡�|����3X9��u�`R��gqyZ�[T0�"y���:S�ȯ͗��S�vj��QLKc��.���V�7d���s���?i��~�m#)�v�y��F�e�-1����';o�Z	��@�=!�n��j�R^�Js���^��a�wY��M��y�Z���J�v���q?���p����&��Q�!�p����~;"����O�q��3��ؖ:��,��[Y��e��� Xh����e�)���a ��:���F#�_څ (W���&��ɔ��x���KS�MG��ͺ����t��N_��ػlFf[<?E5=�A�o��I-#Q>�+�����q���z��Dk]<m���,����rZ�,����1"3�zUp����2 �X������c��B�..i��rhvd��;��*�{�7!�i���Dk�n�8�oՖ�</9V�G/x��c��:��/ƫ��������豊�8�3�@_�%�d�zfc�n��!���@�������at��Z�F?�����ʍ�s��u���Bvi*����W�R<�{�T06wq�E)��8at��,k�B�$H]%����Aթ�����^��g�8�RR^�[PΡ��edc�O�g
sj5��G�m���R<��`?����W=��퍨�w1=kl���m�l�]��͖��k"9�*��{�N Sbː�I4Ei�&��Pdj�u�0EO�!�%���$�W3��h�rE��K�K22�M�DN���9�ЧL_���L�{��K�I.:k�L�k���OE���A'�	]k�A��A�ߊ�|�@qh�j���c�z�ߨ�y���ԆA��o_��+]���2�34�d���E������o�$�qlL_urG�V S��)�͖��n�0yng���e.��WE��7����y�M�J N�P��TX(9�.)��,C�~�u���l�U���8x�''4F������1��WXF4�ҙUⵋ
�����#����p��@�R]�6>�^	qդ׾Kž������h��-2��-/����YjyC�Okg���:�]��\�<�8�@�u���d���qfNw�R�[�fy�ɶ)�U��N~����AH�+(�kwQh)M���i�8E\�e����wO���s��l7���>7tf�@��e��T�
<���K3zt� .�SІ1�$Z�y���O�N���u�iuz�n�dk��+Jz�;��LN���vT��h�Q�!<2
j}���, �&�駦@����zyA�9�m���@��u1��:���Y���d�f���!��y�ݭx��R�*[k,[hm���_�ܝ.�K��麫��$NJ����q*�/;[��	����H��,��"8��+a�"��� �׸	���~gG\��_ܷ�q��P���ô����|]XV�إ^�(�(�@�q�Z�+�!�	��5�S��E�v�`*nW�K��mL�f�s�wπ�=���$V^�k�QGg�R�,��*�K��=IԲ��Ȉ�b��Ȑ �f��6�<a\e��#�U�jiMTI�n����aI�&~-/���g���~Q�b��3
��h��gS{�ѷ||�$zt��>d�$Ɯ�r������}���&n�/]F�f[����A�u�	ġ��(����v(@Ɏ�C�9�Ƌm`��
�.�\�������� 0
G�nѩ��-�vf	�G��S�y9�ƾ���w�L'E�hZ	�+Z��� �U�o�ӟn�*t��\gP^�Ѷ2p%�1�	L�s�|�Yi���u��U�7�c(x���[ H�'h57��`��_N��k9����"}�|!��B�"�����誠����{`w��k���{(�ӊsV���v�v�?p׹��Huv�=p�;㖍��ןP��I�|��!0�������M�t�c� ���N������-��O��8�T�g�W��WA�r3:d �f~��#����*��Ñ!����<�D���V�!��u��+uP�6��|Bd���"xY���p��g��)����!�KA��Dbת�<�;�2�xl]ppD�B���8�W<LD�F.%u�ox�H�s��Ƥ�5�Z��3�v#�R�T����ܘ�sl���{��E]R�݋O���\f�)�%w��$�h'�w")����N�v�����tG��n5OҔ'�\$��!�=A���v<���}���M�k��#�����Y8G�sLx�u��u&u��`���Z��0ɺ*�2J>/H�)�_��P #�XC�<�UN����0��S'�E��c&&KW�8�P�@�Ƞ��}R�56ꞟ�s�򪏶�ar���lL�g=�4���6e]�@`/4��t�]�F�:��cCFD&d���Tc�:Rb��t-���T;���-�#�Nq�'�;�t��T��?�L��M��rbL�~�S�.�#(
����r�^>?�$�I��XC5���>9�l�2�4]�����r�]E*֨X��B!���I<��8�0h�1�{Ͳ�z���Q�=?��|*�����<�^ �yɔ���'jǸ ������D�F�[f*�.��J|���ˆ'-�Րn�?��E��}Z��4h$���j���5M�3��:���^c������ڨV[�Lb?���sě��H�k����	�ب�	�'���WT����￢�H�cX�(������Q�?�Dp4g�%F��6�� l���5�.#��\���tS���ɣ���Bc
��*���R4����c���Ai��sC"u�)s]���%wYO6y4Bۜqg�oŏ�G���ء�-3�����H���3��,!f%���� $�Y]��x�i�*���;��AU�1߀�Bdx�[�����H��v�X�P����C���4n�q`�?70G��ua�Ƽ{6"���Yn_AĲ 8kY�}�8�B����R�!���vj���L{���D���3ȝ
႞x̜�bC�ѵN���*uN_p�Via�����z�ŴY[׼�1�ݴ|j��H"��EE7�a�B��9�㏣��É��������Cl��ǌ��qc�I���=}��Vb���`�@�M�U@2wy�/��D4��.�����@��M����Rw9aøZ��\�BŌ����nb�C�}����=ѯ��%+(ݯ��f�Ibև�%�d⫧�[�=#�[����P���G{S�ހ�$�;:B�8��$����WF��R���z�E�q�����=O��v�R;_�"_�&]� �l��d��w�H�ꨯHY[A�&=����p	!N�� �R��Ɠ�.D�F�+���7�@i%�j;�AP�Ͱ!%��;.XBlӧ|S�؀xK�SRS|��W���w#l�6�d�&����X�ݘ���߷�����Q-<������=d0{���-�5�q�.��n\x��B� �>r�<(�,�1-�IVi�o4">x��{-O� {$�]�.��%>`���_��t�k�8&ő7���Eի8��V��R���"ԻGћ��-�.�%Fҝ������qZ%��Y�S��@���x��?- }Kp�<��	XW��^w6���ɻ#�,�j��	p&�D��?!L�������`.rdڂ�}p�;e�ޡ6��S+�m���8��f~.�QIh\;W@�$+�cjO���7��>3H����d�za��ȽbT�oP%-���Eb�&��Y�j�~6�N� 2��wUd��
�!>	���A�=d�S�[Y��.�}��	�^�of��_WA+�,��������7��Q��:�z��I�Km(�\�2+��ҤU��hԯ#�N��a%�71,�%t&o���RI��ͱ*P� ��u�YH�R��O�u=̓�� }��kmc�ȫ�6�"�IC���e��!�(n2��`֖i�j"ZLR����{�[)�*�P����ͱ�KD_Gkl���Q������b�����>�d~�ݙ�E?M��3_�{Q��VoIB��wP�Bԫύ��΁���߅�1X՞}�n�������%D�n�;r�J=ʁ����sb+�7��H��M��M�ފ�Հ�ؤ:�GF�BEg�)�!�P�/̩�������]՜Gm�4zU���l���D�L) kd�F�8��A�?E�::ph!��aQ��<�4�C�H
���!]!Υpx���K���8f0gT���m�0e�o�
)���Qi�eܳ�L{���v��w.r��J�67e?���&�M�$�rO����||̮�2��T�@L��؟�����v3��b���pzm,%��Xgv��~�p�)Ĕ7LD����k6���&pY���f��]Q�|��v;�l(tȮ���`k������X��R6�׮d��ߦ�H�p9�7ŖX�U�f��I+���<����1#v�1c��5�Nj����n��.c���u�r�;t9���-C˥���qb�b�LYu���~����ܬ���ޭ?}z嶈�E4��=��+B���|z�gg����P�����	�>�b���h4W��=�Nhc�.��MeX1&�:T,K���Ҙ���p/{(�z輅٥��&ܑP�EO�9*1��]w�0�$sG�4ԩm�d@��Q<5{z��ֶ.�+�
���&��@���Uyh����vn4x��&��8\�F���QB������	��P����>���hp��$ ��g�;�9K*�������TJ�9��F��~�cd��;[�}z$�#�u3;��]CZ���)3`��B>�D�w F���������� 8���e�с8�+�n@��$j��T�q���w���D���'0@Wg����9�C�q8�E��Pr��c��|p�\��T�Mg$���R�pEkr)\s%V�P&�f���;h!��Y��<$^֗�(�=���:�#��dչʖh8�C=��F�����<�Ȝ���D"���Ǣc����c��EUXщ��-��+_��Yx�^�M�ٌ?��J���އ�~��y�V3R��`+V5D}j[L3��4�\x��yX���}���Y8��u�T[�6f^kIn�J%^�x�*�j��{�C���ɨ��CEm�s0�K�r�P��o9�֊���>:�Vgy� I��3c�Mp$���9�*-P�8�Oy�b���f�n.&�ӛ�}����W`���c�c�H>^��gP���4}������Tu�Rȹ�1*����������X��bY-����d*����e@7�$E��:��h�G&d�����/'۱�@�����?=�( ��:M͢ �\�o����r��|��Svs��i���{Φ�\|�	��^\޽�+�$;�Ď��Xohah]��s�$��F��A�*���.&�r���62�lV��!�J�J�"ٙ�_} �pT�Gik��y����]ܐ�̟�Y�0��>.��}H�������9V�6���;&�%���~Z�H�g٫�b�@8�v
�\�!�d��S����D��@�x�3���d�Q��W<��YѦb�`�.ݕ��#~�ق���no�����9�Zݤvi�b_���!Z� �&�4�|~�R:M�!ķ���3�l[�P���ͷ]�o�V�̵��q�̓Ea���� ɮ�#�k*P��=� �c��k�_3Xq��2N�a�j�K���Lx�UkQ���\��P�mS��T�C5׀�Z�N�O�;��e��������S��3��~W+�b�t]t]5��I�^�Eo��#ԋ���\�Htk��ޖ�4));-��f�n��������ml�s{$vw�Ei=��So\�ѵ�#�+K��������<Z��S��������4�߇1�)#pic�W�X�`��&	9H��y�//=ӽ#��N$�C�ufBd�ַUʰg�$�(tr>Whbt�a��#�VKohF7-7
�o�k�t����D{
����縻ph �7����e^�t�}ӹ�>�G�㿦��K2z1�g��S<���=�ց!�F��^�ku�
p��D�e{���E����x9�Ս8�7���!���!P[p����n�_���g�SI���rBcx��F_����hd"����%�o0�� e�&�&[��Yw�ĭ�JQ؈�|y���=L/�<��B�)���x�}��>�ȓ���������0��#GU�������<6�̮KE�ٗ/@֧:�81�a���ckLb�˛�j�yI/0�&���r�{�<F�m�ք0M~���*��g�LP[��s	0���d*�0˦nz?d�$2#��8�_�֪���$���a�Ea:��L���G�A��l
��39E󗝛��[uל�|�&H'y�mZX��~�=�S�2+7���d4� $�ݎ��ت��$�2>�a6�+6�S��������_X�p{2�y��3� �3PexQ�"n[�H�����OAE3�8�մd#3RI(����oj:z���g�^������W�
�/��
� �����W���e������
�'$��<�$�-���U�ט$q՟P�!.��Sv��i�/����>�����a�A��9�ơ:2�U�H��d�t���+7@y�I�7��A*r���VRc�XJ`����PK���Wb��SA����yޔA��),;b@�i��2��a�;�.����Z���;�)�';�R<�C�F7���2��F`��)NJ�ه�g`Kb�Ieb~���d�K����J_�clNl���4�)V*�Q!��%H�t�CŶ쒚��O+�Ԑװ�^���hB�2k�~B�Z�ʲ��v��
o<�$D)y�A��ɝ���:g&�vԹ7��6٥ ��w}�ݍ3+�# ����M��6t�g���H��9E��td�4��S�j��z�<=�묢��#`8b�1��v�"��^��m�*��GR��.�Gmn��Y5_�n��q�)6�;V��1vQ�L�v�T���:0@��L��,cI-��CY�bG\�i�d��	����-)i\�~F�G.(�k!��~L؀�\ʋGJ 0�b�GϪ���\�HF�����:C\%�"�>mxm�x�Y6Hç��Q����4پ�������-��ل���xn{�%�N�t l0JTH�94���e�pn�	�Ly_������4�o5/��8�4`��;C�
�	�!�'�IUԄ��v	f�V�;���$�K@�0�F�~l�Ƨ��<Ŋ���hJ�J:�)�a�3���O��^ c�F�&�@<�w���ȏ��+H6X��œ|n��c �����GY��$�Y�%4nLG��2é��)��L��1qdOu����^M�:9�LY��$e��c6k��i��.5I�[�yZ��%A�T�,�Ǜ��qʍ�1� �F����Z�K%�/� �Tߐ��c�[�q��6�w�D�e9������R��D���r58F3��m[�.��^��v�����AT0r�����ƾ�9���i�r,�Ɗ���_��>=1��ug���}��m��CRS����YN��.*��l`���y<��k/F�K���=$�S��y`����&�XC'�:��7�9���=Gy�o�a�"k��<�A�\d�A�[>��^��*E�l7�~ʀ�9!�q.�Oo�B:f���t"�zB��?�3��Q6����F�{πE'j#n`h<(":�gf�nR-�ĉ�[�m��>VP�(羭�k��|`�/��#��� $�j�c�vm���[�S���}Y��`%<��W_,*f�:A�T�+�)J�߮A�9����i��C���d�Jr�l�&ߚ��=N+Qi,�c·:8A���k���#�\�ӓ������Н�3�2�B��j/#Ai�;���@�0�K��cd�bFd�]�,�^�����О�;H��'���Y�S�����>zY'��!'���_E !���������9�s�1`�҂�_4���W�AF��a�9W�P��̀������1^+�=�����"i�Ճ�ܰ����͐d��T�:�XY,a���v�~���f ���s=���n�k��͓�p��B�HU�I�ݥf���Q�<ybS.4�A��/���dih�WF\�>"��S�I�G��Q'�?/?v�,�07ع�nY?���O�w��ު�F�����_�I0(�5���,�����*��Cv�4��(H]����l%��ʹE�Y5��;��]r���
�%l��/3:��q���@�3X��e��9-���ۍ������^>���.B��m������@�%�'���)m�]�敍��5�B.�ތ,��h�����U\jq¿�ы��w8�67��fJH���­�H�󑙔T^�0a�xu�		uLšFV6%�r����}W㠋$`�dtR~&)�����9$� i t1�	��������2�_�����SL]�lh ���ݦ��F�P ��M�����T>U��C�\�?��x�?�,р��@��{��o���	��_a) �db���g�3�T`�Svŵ�:���5/�֨���
ED���'�*PPX�\�ku���R�0gT��a���Կ���,7��Ǹi��km4�@9��m@���$�g�K]�B/(=r9'�œb��`X��j����R��<����4�4�!�]�C��0xh���o;Qf�����ѣ�d�ُ��2��*=YTqj�Kgɸ:C������7$J�]l�sd�k0�t&2���F��mK�2H�����P��v
� ����R?F�5�)�9O4GI5�-K�R��@�Yѻ���dcO� �Ԋ1�X��}��u����8]�.#B�҅�cR�`+��Ƹ?��ǟ���c�u�ķ��Pq���^���w=���Y2���~�c�_�z���Ք �a��:l���]I��m㤴w�+�D�p�
{vW �6~�^���w1,B�Xꐻ#Ah]��	٢.@��&K��<@��w�� =�����L�NԇȬ2�lFΕw�j	}�f5"��ܕrNU�,� ��p�w�֔��T4/_����R�ɗF���-e :D:ON�t���Vhg�-�`J
p�%erof|*c��`Y*u��:@wǝl�e�ǔ��J��(؍��<`%;��	�~|뒴���-�`�`�Zb�(�H1&��u��G,�S�@.��[o۰F�|+����K�V� ��.�Bz��䣾��V��h�e���ʩwFh�Y�i߰����I���9qU�W��~$�����f�I����BCG}].&1�Ի�"qc
�t��0���:$c��*"K�5��'/�q}_Ў 0�zS=\�&�x1"
:"%���X�
�̦I��A�;��� ��䫜���>5�ҡ�P��>[1|e�-<��~d��	�}G*p�m�ky������f���ڍxEG.�\)�G�
QE��;e��uu��2LJd��� ��/Z_��δ*��Ҽ��3���=:��y����Pv)3륶:Z��a�N1ַ�$)�zHLD"W�{����E�tA�W�<�z��R��6�ʈ�"5\�N'F�%�簶I�Gn�����{�=���rZ�FQ�Lc����^L�d�ؕ��/�S�@�|��l�N�� �����1^�Li���3[}o|	�c���Լ�jCur��#�0A�Dp��Ⱥ�v"��gg��7� _��`&�r|���
���l+^�Uȑ�{��9�:�U8%[��d`�L<��b��x�У-���U����*�L}�����������o�N��q��M��m�q�9��Rʩ�L�ʗ�������tq�P�kbd�Ѕf�҂el!f�|s;x���N�gU�� �u�#��7���H/��5ϧ�d�T������~擾{��B*X����e��92������R� 4n���g���M��#Җ'�R3��{�U� 2$?�X��)`B"��RppP1����1J�'��X|��k�y��u�b�Dr�|���*��Fj�0D���j0�7<��Pv�6�e��"@wW�wA�k���Af����[Y:�. �&K�4#����Er�h͜�F�섧�<tovﷂ�/G,B;��Ԉ��� �H�33�s�C~�:l�	YV�����`�N˝��"��eo.L��eE�v��S6������ZŅ��+*��c ��J�����6a��M6)A+S 戤6Wi�$ݨ���嚥~T���(��%Y�զ�D���YX��H��)��>��K-��݇W(Kɔ�jYn=�"0�]��I��;�3������$k��V�/;~Lp���X)�]-;�$E9�G�V���͗hy~o��P��m��%�,]0;���%��hI�R�1���ؑ�@���G/&�$VҰ��Z/���K<[�����%���ƒ���PP���2W������\�%��`�����Y�=蒜4s?(��]�x�ͮ��� ���hK�`����cߟrÃ]r��')�ؕ����*ھ��V5�v��1�`�����)�e?35���,���x�Y�O�ɳ���#{��=Н���Y��N����f��;����S�[V[DHtI��7e����1X�ش�� �4R�N�UFWKe����c�ڒ�ud�aN�=�FDԔ��l<y��o��YW�¬�ܹ���ue�ź������4J���k�O�2���;�����R�G��6�du���L3	S�8'-�AO��j���!c1��Bq�<]髅ü�`�gex<��~�?��oS�C�I}�o�H�o-/�έ�;Q�����~ �4��d��P�{K��'MV�OK�$`��f��4�>��%Qq�Œ$s����;ǣ����<�2{��W��Pl��Wg�!�N{0��w�p[��{���7t^���(M�L�����|{)R}�Y	�1�"�8n����$2�ꑑ\��\�ףx�,��ѩS�����?&X����7�2�Z� �=������}ܝ�ፚ�!����k�gy���O��r���R<�>�iߝ��Ht1p�FLd]�al���c�����NT�bD7���wlЬ��� ����-���c�+��N_{�*�Y�Ǡ,l��]�� �i)jݶ"��~�_<%�q�����J�n-��.@a/7��H��d~(2D���n|�K{]�y�ԍ�$����#��>s~E\@�E�L���[�z�go-�y����B>��!����2C'"�w��K!�@��ANj)�
��B1�R0�*����u��.�Rƾ���/��0���=:�� �$�i�Ⱥ����"�E�$y6�^c�gW�⋙by�O��91E����%�["�}C�<�8Tjv={bm#a��C�ld#��^Μ d�醍ֳ�}e*���E��b�2���������īɋ����;��w�� Eg;�6��v�(�W8S\Cq虚��~��Z4�W����4�-{��~{� �PH����r��J$�4��Nn�.���y�/_Ǜ/@�BR�Rc�����h�G(��$j�&͍g!��`p��#�ad����amm�´��O���z�1�܇��f����2T�.��.ԡ��`���Vǒ�� �ܒ��D���l��g�t��Y%����s�˨ق���f�����$�p�VI+s������3nɒMSp��{�Ϋߗ�¶"kO�)�8�C" �+Dqns��cO)CCb��x��ھ����p<��Z~_�ufi잿���BO�kʇ�'G�J�{ѹ9INAa��k���Sj�=����E�-Q=>o���T����rb]����\c� �Qsk�R�Ō%Q���n@�n`M@��Ƚ����K��&3��l��3z&M>�d7����y�y���(\�T���㒊��X,%�����HT��&#���]�bA�Q��{� (��>f��S���Y1�"j\����W$�+-e�Iz�)D�c�<Do(�TQ�40�t4����KH�Q�y-�	��AT���:�uSC��mH��xp��5����x�(�	�|N��86IE���\!kfǆ���n崡���0��h�ģ��~Jw#R �Vu��A��nZ�܋��t
�}�rX{r!�-���]Zf|&E_4��	rLt�r�.J�ѯ��\Ӆ��w����5E�A�/̠m7=x��m�����>s�΋y�)N�>I0ȴ/��s�u�t��/��5��CwMDQ��.$o��SP5�Q�ω�w��5����}h��[�����>9q�9�9��b�:��$҂@}0��|�V����@юdyZ��j/r~�������֯r��Ft���J�r�5������P\�yʣ���nÏC��]^B*�y�*�q���5܄��s�䊼�ǀtܺ�ϚnKz3�,�?V`�dA����dg	� �V=��wJ�Q6#<���F��K�1	�Tnz<�7v�WE^s�װ�6��!�]8p͓�M�N��v3C�)����Fĵ�
CR��G+�����q���C�s��tpA�O��{���P��R4��R{URZ��K4�W���vu������Vs@�hv	rQ�9G!`b�Id�8_��<�^hfp�
	jy{Xb2���Q�-�5��Loݤ�k��خ�6�J�rH��"��bY�Zq���~p �1K�8 w�W�xϘ���u�x�;�I���b9~s�3� �lӁI �"d�Q��Wp���k�sK�"*Z�9$�C�jG�b��B���b���i�ˡC�"m��tG�z�Tl����)K���t$q��1�1;f�WbGɊ�Q>��A� O�x"ª�Oc�Ds������p�qr*�9k��2����l��c+� $�SYe��.�[om`W�s���+}�����j�9�(}�lz�=p�hM���|A�)�c@,��V�~���XG��ĭѢ��@jN����R踇o�dIsWD�VmcЅ�BN�L�S��G�\���1)�%�h8Uy<�
�M��,�6���Ad�)��5q`�6Lͮ?ݱW^Пf�om�1�f������<�:6���z����[��Ÿ�z>[K�H~MQE��9�q�/rM�x�-����u�`���{���5�{�͖ٚD�/mr#�$����R�ӧ�߁��EP�*����c�kSɐ*��M��� `۞�ۥդ�o�p�gY�ƴ���pnɢo��o\E����@1���J��7} ��
�}J9J�'�n�և-��y�#�)H%�w;��֓w�����G��G�1YT�
w��9v�H��e���ݺ1U�#%�G���a�\����Bq�$i_v��b����@��Re]����y�!]��YvK�o���`c2̏M�;ꡫ�Е�����)��7E��yk�d���tO�^���u��X5���88��^�7��ʂ�4�ْ�zm��숂���.�Lm�.�����yƧ�d{��X7j1�T(����TK���v|�EPFW�J^�����v�p��#~�΅=.Gm�\��x��z�Y~�BXb�Ә�Hp�M�y�`)��YY%��U�˥+�ŭ�,!�?eȁ�k���T߂u�S��cP�����P
�����U��J5U��^���C�Я����1,�#sM9���&��-1�l�o��^�H���f.F,y�~�X�:�T�������&�����0j��k�U{l��\:&��x��N�r��4�ق;��ꍀj�>fk�t�»��ɂ6���d�Y4�LɆ�SN��ǡc��ԅ0&�HD*lm����F�9��߶]���i&�\ń����n���z�Ry����-�\mZ	~��n%(W[4C�I��OI��:�V�o���$^DoZ2=���ւOB���cT�f��$<�A��1��� ���NG��-�����}'u��K#�Jz�m��Q)�c��`��ee����f;������)�3|�i��n߬
 �R��D2�W��,�7#�c�v�,}�#��xҊz��E5c�l�"`oez�zכ��&��#��*^��a�`�v�%x&J�Kh����z�Xlf�3�S�oT'�#���ڿ��9�,��%N|� [╆��-�Z=!�o2��ٛ�o��@a�^����HFx���Z��!)R����(7i�̘m�/ݸ7�io�.?k�O7i�����29�1ciY�mLʛ��&f�C�hI̘|��ҵ��ɧ����{6Y�>�����´�!�C�6��^�y�o�R+1"��θ�W]u4Ʉ�xQ��'ȭ�	w��%�
�k����o%>D_��l'�WTH���nGHQ�^V�%h�t�<fwvj�J0�)��Wð�Mq�3a���p��v����u6�y#c}?� ����(1�Q�q>�&�<��Z� �E��%@4r7>��4�q8?�A�����������yL���4��Y���>=Ʀ����Y�T|	�߲o���i�������9_=aAb|o&�*�,O�T�w4~�MJ��.������b8��ڶY�V6��U�q,V�W�mQ�4a���>���l�D>�|�'�	��d�_v�x���:��l�9)�b W�'s2�Q|�wMa@�D�i�_^tޡ���">����(9ů�'�1Q?B Na���MLq���xP�O���t�I�Vu˳��b��@�6�P�;}�3H��T��a{c玮�4��D�7�W��Fk�ܖ�!E�渴�������~��`
�3
W�8\��[�Z��Z"�4�{.=��eq�Q��泓�+��Zk�lƈ�����*���/���n�nY���X���Hԕ}ڍ��t��Z��1ڍ���o��������1�t����E�FG������Eq9�=��+v�q_K@兗���
��Й���9/DV��z�� �i�u�J���ojI"x��d�� ��]v	r/��LѴ!n�~/`ՒgO�ʩ��9�������~U~K�YJ����Z����k���|�a�.� C�,��>#��z��OKJ�g���	!%4�٧\p����y0�ɹ2�q�<���:��U���dq �f,eF����$����09�L#��oҋ0֡�ӏ\���"�ꭃ�6���(�LaтV�1ڿ�q�.�΋|�!�}#A�a�;�X;�;�O:W���Wmg��(�%,܋8�������6yZ^��p�� �)C�R��QH�1^���U�hB�L���j�l��v�ٝ_�iǇPt%,�U�N�`ب�<�u���#�9}�U�����,�������0�.'~I����~�/s}�(���*�-�ϱ�4ֽGd���&�C�� `@R�)��
p5��e+Vz,���Ǚ��ʊ�|�v�KD) ��-b��-���<Yj�0)ض��v����8e�9\�����qC�+fi+��ل$q��)�����)>�Q�)�?��GZ-��9׼Q�\-&�BJ-̖�4%����D�?¢a|<���D������sT�K�?'�mL��.�C2Z�|�|����
�6��YΪ�������ފ;uX(sF��>#~�K��NoqE���+������JyYص��m5��jeM��W��u�e%/���^��2���"y�̄;�ےQ���S�5���m1��[	{�0ʼ�h�|�LQ��Q�� I��ft}�t���>:˳�Un�x'ɻ:���&EA3"?��w��?Li�9X�n�{��P"��d�{�%I4n�l����z}ռ�°����1+���ck��X�w��&-4H K4m{̤`�����Ʌ�ެ�i�g+��amq�跛?��7�1�D�#)�\f���1z���#�s�qy�����~Z����׎�i��a#��}[a �WfEdrr�OqnB�J���K2l��!�ݣw��^��{�5��=���g��jO_�	u�(�-�}:�8z}���$;S��_Z����3.����D�h�]W���</�3�Z� �*��%��_\��q�&2\͙͈,�4ZS�Ů�3�����"�b��l�8�����*��e
G["U�c��
�-G$�*��4����[S��z��*�B�x��W4�{��%�b�?���(�EX�l}�Vx��g���1��.�iwo�5Q���2/��PФ)��e�5�Ys�ۓx;�x�t+o� �Oo��N�'E�~q����-����ج:�z�ά�����<m�Н��d�7p^��h"��)}��y9R��޽[�n�t�B�7�7%�� �l'X?^�0A�-���܎�h�e�3�g�t�CQ�	�ؑ8{�ujV���N>��x�^ɉ�U/^i��Wc��dB��]��V0H�����Eg#'��Su��[�Yd������|�j��)ز���v3F�Bp�pL�>���_b]���8���]ۂg�J�x0=FK��)�kBд�{�:�$����n����D�d��E+�3�ea��"�k5�`�DH�e�K��������eK�%:{��+�IǆnK��{%�)4��K�"s�Oc��������̝�0���[��{z�v��`�Q��o��]bƜtZ� ��:w���ԺV�,
y�*�w��v�G���\kdN�#*o�IY(1]�h��=:�0��`hБU�r�k��~�E@dyL���&AbIu)՜J�(X�cx���wA�!Ӧ3��t�m(ɠB(� tl����m�m��[���z��'��;��f�N&t�T�W%2�Jn@��2O��1m_��_I�_���W(���m�V�F���U��Dy�x��zb�^* �&}��L�Y!`�fCH�Ң3��M��}6�v�_T�*�CF��^����d	�]�L@�U����,o���}�A�!U�\��r�"�M�v&�9�1!�bPt����b���94��H��Ñ�`r��F���T��&D���{�k�#q;XU�2{���M��0�r��ߋ���:覧�bI�_�սs1~��Z��}h �f^����	�[8+��$yqճ�e����G'��q0Ho��J�Xʅ���_��lB�`��Ka�s -g�ߓ��S̕=9�i���v�j�C�D�QTĚz�T]11W.�_c5k��h�G���ｱ��ڼ;v�w�x��0���$.��&ꧬ*
r<9I�T�^���8ɺw�,JuM�2�.�;�u�Ds��r(���Ò[\���B����Y�vO���loD#�ck���"#�h��.y��r.S������Vq�>���������	� ���_*R0y7�8؛S����q)g?t��m!-�o���]mcL�6	K�A��(�
�룢~���Ё���8I �u�ˢu��Q�u�2I�T*��@E��+�ްr����բ�.�3�H�}^�L�#��!{�"�=�w����,C3�9�bnG/�򮥸�W����z庨s�1׀W��b���
���4��A��H�Λ7
��[ޅ�6I�tG��e�����~:M�m� ��yLE���,x��Z:i1Z���mif⭽����3��:˹�7��q�c�4��_nA9�ܼM_�NA��wM������Y����[�F�i
��H�{�X�ИP�=O�B��\�PS'�`*�݉���u/�lԖ$,��k�֬`e��V�_8��/	{��
3씨��S��%ϟ�?��ɟsM���|S�A7�Ue��P�i�s)��ٟ�7�]ǒ筘�3+��W#��<�j���
\��|3?��oέ �k§��a��}�)�fJ����q��^�*%�L$�~?�߅9xF�tz%;?���6���ړ���������HzN���)�D��T�ׇ0��.! +z�	�=��OӾ�*�L��0�o�>I���/�σy� `R���1��6�42���VБɫ�Ӻd�Up�h�T�׌e��ݙ��Nl4�i���7��^����p'�����M̏�'�H��E�J��mD-G�A��#�"��瓼���8̲�@o�@���w����ӆo�dUn�x1��&�U�e��jD��+�����P��i[,}�S��yo�6�� �@\h��4Q�0G��ĸ`V����f9��5�WQ��]wʁ��A���]�Љ%�-�̙4����:ܲڐ���0�Kb��F�Ǝ�C\�8;�ir�7��"P�)�0�g	8�FD�^��޺v�VW?���P)����P7����e�DEf��a/��(y�1�I
(s�Ƚ1y,mhŘ4bJK���AWO�B�Ǫ8��77�v{o�T�,_���;¡�;��fư���YS����+kzj�9���㴰S�V&P�*���)�K��k;U��yF0Z�4̵Hc�ށ���(k`�>OJ�o_IbM&l�f �c�\{�1��ƅ�2�Q�|�bw���y0q��~K�����ef��J=�V�Deɝ:^W3���l�Z�}2�����=K�� �*�j���3�Z�����7�$w���7�eX?~ e��Ye3��MK�Y�z4�K 9�)*C2�oV�P�a2@^2 ���f۰=�B�p�J.��rcA2�o�.��w�:��4�8T�˯q^0����M=�)��VD�W~Ρ�~�?]�K)�lw[��0f"@Ԯ5WZR���qz��,������0��0�5N�n�Y�Sӊ�fO��)y_��U3�XǊ�=&�d��W{UBXI�~4	�k�U��!�8b�����H�5��c&)`��E�5���Vuc��\ƝƝZ��^�vb�ˌ�z�v��u��f4D6p��t�#̆DS�#:��;r�a
-����At�*�y� �:M{�H�k��G�[$z^2[��ʪ΂N���V ����W�M���q�_���<-��o��o��;��g��t�f��f�D��@-��D?5)�F�6�s2��T�1�����?K�4��UA�
��4��eʖ-�N��M�ˡ�]�W����u����+J�s�,sXB�����6�c�B�$<a�0EJw�T���SцX*���;fX�ys�bP	�l�ՉQ�OE��`��*�|�v�53��%_����fHּ�}֣x�.	�kYs�&\���� "Zۍb�W+�틄mc�IՇ4�^]�� k$áu���к�w��l{��L�/�V���i8c�A�R3�=�Z�R��E�6g�<r-�[F�2��4�X��<�.�G��d(pu�:O�{�@�ʦ�2�\�&|Ruڧ�D"�kx�%k���u!N��E��yp9(3�ߧq>�	��e|BW0t�)_�$��؃�(�d�3��Y�#p[�p<Q�S��p�R��^��X�pa��\�!E�U��R���X|���'��#O#��x�T�x�����oXR��ʄ�a"���l��l��K���^v%�J�T���
�о�0ๆ����`Ea ��(�$��L��wΧ]�.K��m�m>�Ս���[7��%�2#-_6x��~�K*]�o��Q��w�u��Hˢ�|65������l{��$��#�����pXKƾ�dJYr�J
��`��b���$��E��j�}�?<i:>�貛w�U�T8o�a~���;	:D��a��vW��n����*S֤�;%:)�;��U/�ʄ�PG�ZG%2�5�}* \+�g����鹪�Cչ�M$��]n��]�#wX(;�m\%�L����c���V����UoZ� ��R8�Q@�n	�9��yH�O-´�c��W�٥��:�:[�6�X�ZC��r�(�ܾ�$Qzwt�}~!��a��@)HοI��I�OF�����T�[�l2���i`/�p!�,��ޑ��:�
6���)���-m�'sJP��)�����	V�tGXt�W�Ϩ`�����SWz�OC�[�� ,���.i�Z�'��_�p��\�I��c��ʉܠ�`=�FҞ�N� 2��ޡ�n�_/ZR���(u�M�lM1�m�-Ԕ;����1�-��B8���� �y�;��H{��Dt�^cl�ߖ��F��S�$+�[�f`�v<�P&_/���XK�=�Ʊ�7|����/He���� $^v%aԀ�����℈*��r�³¹��x���rL���\wMt�3�K+?�ء�;2)�B���C��O��"�0�-Z�!�D	�D�N��/����+���v�o%\����'�$S���
Ԉ�����P�M�����IaJ`E��t?��������l�������آ���d ��wŢA�üԃ���1Ad(���Ζl.&�c���)�������_W'hmRz��T#N����1�������,��.H;H��.�D�G�	t����`���O'��:�[Qe�%�Tz~�X�hN��uy!���iv���������s�<��u�v��X�kxQP��q=T���?��X�S�?|r�ͭj��=H_��:ku����vK�&1��m�.Rt�m=�ѵ�ڳD<;�:1�q��v� ���]��[�MBГ�6K��ǂ�i��A^��o��j
��@���,��
V�q��=$�ݤ8exUe`�\��-�����x����W�>������2��R��D\�]��Q�ni��B���2��?6���dX���I\7a5�7����C���L6��Y�pw�i�r�60	�l BNY���T�,�4>�n�X�)5����&xM�ݥjʺ��*�d>�oxc4���>�������>�L纞<;������;�?k�jno�%(��t��Nd��;��Ww���K���B8�hSj��m�!j^�;]�Z�`fFE�U8�&�WD��P����bf�ݺH=s�4��V���zc`C����)'�
����f��*Z!(��D��}�Q�D��|B�")���*�:4��K�%�@(y�E;O�_�ot�S،�r5+Ì�W.�sq���}LN�gn�aЈ���=sL�p,�����5�ɀj�6{�Tͤn�E8	 �4��+��nH���-�n�W̷ﻡ����z����P�`Ѵi3��t�)�rp�uqU��)�I0_V*�����a1����\����I����_µ�,�%�u�o)%��c�ڴ߲��'	��p�ߝ$6��֑�J��An��w�^���%ѿ�d�� �Ւ��T"8Jm�����SS?�;�Xԋ�tR4��.B�K����}_�������>8B�f�ѿ�p�k�����67�UX�jY/U�;�T ,����=&���Cֽ�B�1��RL��G�lo9��.�q��
P�Df�9�I���"�
6�dsq�V(�����x�B�~�������M҂���6��W$_��d/�X�0�&�4�u,ư1VQ��8ǵ)`�!n�ޛ#��߇!��z����Y<a�c��~ލdzz�:Z��'-L~w�E:�D�1^Gk�y�d];�%���0�}>_���DX�=�=���!S#`�Z���A]�pga�z�Ut��j⠢���uJ-���pXjm��?��V��4A����s_o��zR��P�)�5�T��[��*�~�W��K��;�~d��C�?U�yE�3�ǷEIr���o�W���Z?%-ќ�fP+a�tu7�Gf:AIBpK��2;�`�.�O?E�x��FlqQ��Jyaq.���	h���*��X��<\���h��5��$c̞�~�`p��EB�1B�B����c�NH���UQ���Ttǻ��B)��i|�S��k�̾
<�$!5)�j��m3��O^�d�Qr��b ���C��,k�����\[x�ޓ� P���L���0�ſ+�~���?A�ڳ#g����Y�$�� 3�z�" ��jq&�j!U�VH�!�	�Sϒ�"`�v�0�ȣ��䳃ڈ�mс��A)9�IZ�P���_�^��(�(>��3v��\��l��4���p��tN��{|��x<��:Z���L�x���̌�!��@���$L��hV����R<�K�Ri�Ɉ�[gWC��;e�Y6�0|4c����[)-l���G�- ��e����5�P�l�8� Gh����v8ks�]����b�Z �z̫V`ElrҘ����r�G͌�^�2Ƽ������.T���x}8�D{|m0���C��>�߃��������A�I�f�����g^�h�3;�G���`,���W{���D��
�>��YZzMX
F��[�@9Vz�j�R�'"oЕ�h�1�b�RQ��j���Vʱ���*�ǎH�y���X
Bn��wZ�=C	��n��(?4����iՙZ�[A>���<\H0s�P��G�D7���Wl��,��^"u�"0���zg����ĉr┍�K{�x�9#y�"���tX��i�	��_w�7������a?�l�oU�r�-�F���	��s�e���Z�$�^O�l��z��!�cx�]:⚓
ƛ�;�M|J��-��{J}%��2 ���c[4K�@b}aP�Ҏ^�6H��8h�B� ;X��[����;l[,S�n����H$%F���I*!=����XW��k�#W]>��]W���cq�L���;��[��}��Qu'����vI/���*����
+���4u9���Sb��vL
Q�A�˹��0���/J'��жz��B��ܮ ��n�e��ʤ��!TA<>�2���'�;�%.zyB�<���Ў��=�Ü���@���)G�!^b��@�/�H�,�b�$'���K[⒧��e�]6�-�	0�Q� ���G
�.�W��uI:��ŷ��L����,6��ǘQ��mm�Y��c��M�g�f]����N��o ��û*��(_j�7J��e�He���\�xT���zKsW�%(�,��t�l��
VU����m�e�1�fl@���=���S E�2��~l(��X|D���)��Y�䣏���1�� 4�u��D+�&{۴j*��U�h�����'����4_#j�U(��n��1Z?Z]�Qb��QC|��J���(�^+�6�V&�+_q?l�UҦ2T��n�g7�������?=	o@����<�)���"Ib�-��-D�G��*�c@R�<���n��Mn�?�����u�C_��[���?M�]�тvam�_�XwW"�� �+��g���_���E�ż-�3����Q.���ΊC�f�g��^n������[���3�Aǁ"�_�`����
���<kq��VWQ�'f��-�F&� QPY��;G��4E	�]��F���z�s&K�r�����U)a�(���9����ۗc6���m�9�_/~��GX������#�wF���[V��&m|%�!�>�	���_���z_O�x�*-�f�[e�:K<��.�ЀL���zp	�w.VE*;M����8��gk��1��"AwS�\3����%$p�Q���g����-g<�h��<ei��������HR&�� ��RxȻ���	
���������*�˾����$ot9���Ju�nUg,��`�vB���u)^��a�v�9�ᬌ�k�gźDH{�'|�	䑙F.,:Ϩ�Aoke7:Ŝb��}"�$yhj?�c��=ѐ���,:v�[�\SC|���U峾�=����"j��
�4�-V�*byMԇ���(ٲ��v�(�m�#�,X5	*��*� �,,��X�|��UyD�	.��¯l��e���w����c��<r������F�	d�u�G��X<��T�\�\:i��u�_�#��~���G�N�/���P7�-��BZ(�����10X�ф<ˋ�!��U��������i0ؚ��x�o�����ѵQs|.쯖��
����#�z���w4$o�4����O��N�@|2�0�^���;Wa�覨��	lI��t��ҙȑn��0n�L�"�n�g������g�Iuw�s��{F^��[aF+�:;��{e��x�r������>��22�aH�s�t�#�F$l'�d*V<��d�3�_������	�y?�z�v��ݳ�0�h�������}�����׶�WB���� g r	5��۟��B����4Oc��:������a, ��v�zi��L� �p"L�;lZ�%4��E�˄��l���η�o�?Q�����!#���R'���Mc�Q+!�(E4���Y�	f&(�͆v(0ȇ�D����I�
9-�Lq�ϣ]���85����#�9�i�g���g;��2M�d|��#��X���D-ک�aX�*��Y��Κ2|��l�y�ֽf����\_g3�E���ߊJ%!+�"5�o]���)�����DZ$�p�twQ/��-�s)��H�L�� �:&��MH��n���Iz��������w���V�<撫��aG�QJUL���K������n�Q�{���`9��M�J����R�G��]p����4:��:��L��C��` ����-�Q�
�6��P�e?�^�W8	|&rx��I�]q�w��Uc���v��6��~�U���ii������C��(wX�FV��ͱ9�ݗ�O�u	G�'�)����ҥw���	2m@�GWŇ�3@�}��๭�B�vh>��������(3��g2��*l����bl^���f��Z�Ŭ0���a��Q�?S�������R������$We�̮��V�"ft�OX��4/�KŶ������j�5F������Y������C\R�^�;���Q%_�+h|5Z;���^^,�ڦ�X�i���-�7��i�l<ݤ�Y�!���.��7!�r��rr���KD� ,O�k�^���F]?��a�!�־Ж�|wC�"��>�O��KwX��z`�UgAa�h/k�˵2�}*?o\.	2<`��Q8�?=d�vQ��1�Y�P�>�OŤ$�\��
���|����Z9OW�mc��G˹ ����m�H��^ט�`꺆�r���L��C����3��j�Yn��i%+�Y�7Yy����S��+a�㰗���%Ə,�C��q�VC6�'���Ȁȑ�Q�����+�MZ����L0���o��U�k�\�%3��7�!��Wx�hK6h���~�2�(A8Eۣ��n_�?+i��&�t�@��w���ܛ�����(^�"!�=te��tB"Z�3������柵_�)�����Ƅ(i���?k��C��9���9�c�0P�8��
XY�}^�2�_�\3OH��-ňm��6@5�W�5P��F�_)�#����ٺ��385,�~F���r��i�O���VR#������.��̚�4���>z��v�����g��:|�VX�7���iY��0V��(E�M��%Y��	i�/���aP��=ƿ���z�e�~���*C(��G��5&����ǳ檄(��Z����&����H�A`g}�&�K-\�%�~G�]:�@a<pM�V#��4�,�j!s���~4�<S���6[�|�QXR��/}�����! �;T��e���Yv�2��%�%6nn^�	�˷�Li�C=�p��d�YX���l�}HL�DQ���qL3U�(��_����� -z��.Dя�7���fJ�Y-�A�=�Zu�_b�Ϡ��PEg<���w��XV��նJ<m�y�	��2���VU�De*������U).���Cn!?d3�]��]�w�~.#D.�#� �v�W7����G'�6)�[k�51��QOZV�ɲD׵b燏�,�{�ֺC6�_`���/3����&�#(O�P�d��=x7��/��Б���C-����UX"�U�+��՜
�"D1 ��9��Co|��Z#Ѭ�NTS`�"M�⤀*P/�5��e�h*�8�|��بR�?��-ڹ;�j�q���n����;B>Rd��8a���˴JR�j��0�aǷ>�Z�G�=�� �?��	�he7'���Lf�����P�oe���)8��ĉ����W V��U*Ef��s<���2S��Ï�({T�Fu��+I��Ʈ��(�H��>�;�.��y޾h�A	޿�vTF�Rr��{��n(L��z������Wvvc��sG��P�9��L��,0i1{ػ&ksR?J�x������a_>hN��Y�z-�'l���
!��	G�����$���⓮�/^���绪 ��]�N%�7����yq�"F��*��Y�4��f1�"0�x��Ex\��wuq�2��X�+�����wNZ�[%����a3]�j$����|.���(�T�g͠�s-�E%�8 F5VC#���?�תRZ#��F@����L��C螔r���9[���*	y!��T�C5	���+?�[�B閮[;�O*�;CM�n*�����o�
�7hp���bӑc;ge����G�?�7+x��NMN ��	<��00�F�t�`��'鏯�>	��y:HMٛhR/Q���7��Q���>���:b���"2�;??�.�A���cލ�Հ�vh=m-��'�~\�E궃�P�M��B������p����+h��w�����W��>`��w�ڠ�Ue�-a!f�9�w�\���(�I��l{jq�Jj)��h��,o�޳{j�]E-��}\᐀QC䧵T��g��P�yW7Ƃ
h��B����#~�.1���a 5��q1��Ł`��F{	/��$q�0w����ź��A���8þM�6&r�C~��-$���e��<ᗻ��"{�y�G����}_4WgҚ�@�B�G�}�Lu�D�$5����mf|�����r.1�э'����t�U*B�CK�'��L�^��*7ˆ�2=lP����Tq�)��/��$��5Vk���E�y�K��d<���2�ۅ����$�{bC�uG��c�`�В�iO����'���3�B|�VMi
ۚ�כBDu��������7��AgpxX�}���}�khB�����(^���=t\c���f��EE��c�{�l�j{i�xB�mp�Ђ�k��#����pg��Ś!x�իmiM˥4��&GnRv+	5����8Y��ۅ�����ȭ�x���5~�ڂS�J��O�4ECv4�D�"̶��5)ߏ�c�H��u���҇�̠���~��G�9�ө�om�2ץq�[{�������h(�qM�~j�:�[s����1ӈD�р?aV�@ 
(��=uĔou9��R�$s�i6򻸻Yh=���瞼lj������W����=�r�Q�����?3N��h�*W��#�OW�8e�eEn
q����$�
P���c�cD�Ձz�2vr�>�R�K���?&��0���z��b1~�4��n0���J;YG��Vg������>�4�/#�����
��S����n��u�6�Gg�!5R���P��}<�υ���:48�4���DQWdK*��ڕ�A��44f$/�B7�{o[6J�}i}���G;�4]�kkZD�!���*2����G��	���K�\i-�/Jv� ���}D����`���+�4�q����v��b'q+c���Ie��g-����N J!lo�rt���	_�ɴ�l[��qS_a� t�g����I��1r2��N�ij0Am�;�"�)�|=8^7�Mlnm��nQl�C���X��Xǝ�gr�����St�/C!�3��9șhܥ,ޑWi�"�2�M��Q�Z{L����AO�0��g�,E�a;vBƚ�g�f"�	TW�J~,�	z
�3@����8��X��e�������w���2�v��
�����p�u�R������xPD<h�32�p�e���m�9�0��5ջ�~+�=�J��=ʩ�����&NqL�]+*��(�i8�E�g�\�g��Y.y(�r�s�J0!,��zT�	�֚�п���8�y�PJP*�YǸ�V�Y���N�)�7'�݃W��4���H���6�dC%s�^�OQ�3�6E�C����i#~��3g�00�l�����͡JJ`ʎ2���k�HЙ��>]8�w#2���Q�	NrF�L6�����D����{|Cǻ�i1������Yӆ5
-���PŢ��&��Мf[�J�e=pXS���GG"q��R0�cYo(��xR!Gga�uj<�gx�h��`�d_�z_�d�C5{R�D��DR�1�H�pv�o��Hx�(a#߮��Bhj��8�d<܇�%���ڐ"����SJ����ac���xRx��ӕL�nA��U��Z�ڂ�m��K.�b�U�pz��d�b�|��g�(�?E�����
F��j�������b��Z4��d&�<?W5Y��n�Bs�+�k^�F6F�)�ޝ��旪���(���`'�ު�C���"� [�*($Q�"��C
8zAO���-�1���WV>��e��O��@���^y#�X�O����Fp��w�6�7fr3 ���
����e�l���Y����f�̷���8�l1��$�q?UI������ó�t�C@��G{5'�!J�J��g�y�Ī�D
c*�K���=,�<S��╨��K����x���G@�I�[��t��
u�!��/�=v8��	�3v��P�~�9�Q8	L�`OKXN��w�y�ޛMg���u�]��S"�]�-P[�M}9���2$jx%U�E��4~d��G�	fY@1���_�9A#�̳E���C5��F�qTp�
�|r���Q�2K}�����M$�����A��֖G,��]�g?��X�:��U�F\+@�>z]�S����� ��kFq�.s2����su���I��J22�kq�����y)i�� ��,�O=k�$�����Ek)�}�NΉ��O�=9��c�.n:k�$)?�]�x�_PZ���_����*\��l1lQ�/Ŷ���+yW��+2)N��s�5rb����"��,��ڳ¢��=�/�ɋyO�D��r�7�p���Ywa}�
��Ԓ&��/���J��0��N�+�]ZSŎ:e�C�Тz�e�X�c%�K�����3����^�&i2�e��A<��tXqP5�2�זG������Ώ�&�D7g�^_^;�$��syDY~�}c��{�in���x4�Y�7׳Ύ �WC�kuG����zc��'�ߏǫ>���,M��{�d�N~j�gFF�l "B4�P��vG���Zp�)ӳ�b��w�V�喜�a�K��.w���@d���2]���׳[I9Pi�f:���)��O$�;3�8�KH0}�_#<T������~�@�� vy-�����A��Tl�C���m}�u��X1P�W^ +� ��7�s���ԣ䦕�
���p�}0P�6o�������\m/CF~��d�3�P��%n�L�����=c�'���zQ)����Ӝ}l`�*3�'�G�9:�|�o���s�V��S�q)�:��8_���\=�lV����/	�.,���l��`��,(m�J:�mgwN���h֋����*�ˌLd0�=*�l)���Α�����K��W�j����Tw�%	i�o��,��xE��jSx�I��`'__�N#4\�9���nnY���?���UY�'H<;�):��IB

l"_�N�3�s)�D<s����.tN%h@�3�$!�ʔ�8��lc'����Q��ɂYf��,Dæ?&kb�v&A'A|�Ia7}%�_h݃�vU�T$�����tS�	d|��-W�������P__V����l��-��й�c/�'|��(\t緕�������5��1�xK��u�1�?����Aj�mȿlnf�؊��Q6�:$��~�( Tno��3T$ވL�7�	%Қ}�~���x��~�%!�p� �C������uY�('�e�D�j��������I>�A
��Ka0
(�q\a��}���Y>�x����T
L�ǜ�0f<m�Um�y����z�E����G�����c���Eu|��&�wU`[g��T��#�)��<Б��������t^������A؇O���HUn}�������0|��B�Y=Ҳ��,��>��VE��M0��"�RHK���Ł{]���%�n�"of%�#?\<Tsw&3�r��X�m��A�oǇ��hK�.!e�
⛙�"B��.�q�4���Cf�D�� 	 u,����Bk}�������ͬI^�Q��n��'�t��N�;2������*u�<�>#=*�jk��S�瘞�d�U�? KYr��mK�@��
�FBh����ѢбBf���\%���1�'���Ҏc��-���[�4�������+�6_�&���}gau��<F��i.d�a�;��,��o5F���N����:X������jf�^7m	j�����H[�bxQ�6KǞ�w�@р,5�+��^+�(��`Q����)B䅬l^eNU�Z�CR�����*.�]V���dwr؜�z;HwsŨ���k�����^�Mם�&d����4�9��GG�����k����>�����e(�p� ����| ���OEc;�_��^R�<%���!(��2��B�9<6<Á�uZߥ���8��USc28����۸r!7���;F��r^%��=k����HI@���t��1[#Թ=��/��/J��T-f������A�}syhC($$[�5�3�{(Ol'R]�U$�xe$��[۽�)�?SaJ@Ў�E�U~&g��|�� :���d��)Di	� ��O�]Hr \��q�!��R�U1��s��?e1$[\���� �.W�ě��'r�*�H2F�I:�EkƸ��맹 �"�V!�Z{-�4҇��a�l֭��%�,!�C{���������}��oyȐt�G&mxմ�F=��+�N�+I��E"�Cf3� j&�`gpp:�4���� ԋWg���B�U�qۗ�J����=�~xb��sO��Qh�dEgL`T0l�fY`\�n����_�r���{�X����`;��)�D�F8&�L@�8�ٖu�5��F����̀D�8)���}m�L��q/i.�����+��2�'�=,�]b�Mu�$��.�q,%����z|r���Hx]��M}i��~������77�99���MȆk�,� ��t�If�jG�bvvu�OI ��y��щ�n�i�5��]�'�X~R�!Y��|�jY�@��u�|;H 3f����(�s b�;�*a�xc�/k���l�
kҙQ��`߆�"�P*,,7
�!p�ʈ+��s�S1��-��l4Y��U Q���{��,o��;ֲ�� �_R�i������wB�7�Ǐ�S����5��UW'���ϕ�������Z�kϴ�ڗ�\���I�9/ bQ"�O��/t>�V&�=N��S��8Uk����<�D����Zw˄N�?zz�q��4�6�	Y�
���G��9����*��l����y�t��cJqV�[�|hL��M�bd�g�2/�U��=�#�) 1��k��@�Y&5�m���!.:��R���U?�p�ތ�BKVv[	.�WZŖ���U 
#����N]Z4�f��x��;q�?����3"%�W��b@��"�N��y���9�O�~_��:�|@M�I�ng%?����~��Q3���w�8�TYuո���^��g��g����`��݉�o3*�F5��h>�4�X������Z��2�8�!���Y}�%���8�k'��ݿ ��H+�'ϛ����ӛ�}���+����U�d	a+?����c��B4XJ�c��Aӥ���B+WB:��c��OX0����y��K;+�դ��5؋�
d�o�kjگΊa�LK�ͫ08LN�,&�I#n{�No�io���e�b�)��ĕ-�I���s�$��U��Q��8t� ��Ҿ��ƴ	<��aIdu}H&JE��K2�I�A�D�t\j%��w5�,����˗
L:�$f���Ql�>�,��yQ��R�er"Ώ8"`�K�Л�܋?�'��P��U�������$xo�'��>��pL��]+&��	!����_!�h{��ZH����� I��Q����f��x�>��W_u܍��� �1��X�MS�0#���x�p9�y�"��
}ȿ�p�4�p��f	B�hrry�&�(�|���$���R�C2"e��k���v��	��
C��o?�Kqlu(n
�Y��J@|�cq�qfȌ�w02��{%��6i���Y�.�C�B�G�˓|�@}�n���#|=�t^ݎ���-b�w��_*�Imp2Ĥ����r(���M=<���k�v�/�͙��n��h}|Z+0'@���3k��P e8��CE�b��Pv'���X=�[���4�r�"��Tř�G(�
�����䵆3��T&o5�PO0�p�����x�j��⍸���bM��"���w^4��ڰP�r_��<��.��͟��1B?�%��֛Ǘ�b!�c��U�E��U$i���m����&�鑢"��u/�KY���k&��I�.
,��i5k3�%r!8��O�	6R�&�|5�Ur���oqw+����-D�P�#K��aqf��h7��i�Y� �wD�q��~M�z!����ΫН�m�3߰�D+�{�?�t�A�t�/R�6&�s��+�������S�w��U�2�ĊC�D�yy�ҿ�"�d�N��6r����|ueD�� U���皤���7q�@�aL�-�b�y{@��噫�:_w�5e�6h �b!De�uNg"�V0�C�f28�]H��Lj3��OóIvozE2�A�^�:޿\|u�39�qڬP&ZD'�+e���|�QB*�����)�W
�*k�"��ZC�ޱ�;2�ɥ�i��g?��P=����C�Rj�5X �n6�/���B_5����=G�ۘ�_��.@�����sN'E��Y-T��`V]�!�Eѭ��������3Nh��V����W9�L�����ɌI,���F¤���B�Q-GQ�N�o�݀.����04���l��ބg��� Ti��:,=�p
.��/�����PR.���M�e��D���b�Yz��S�A\έ�\9��ݶ��t��{�w�C�2y+M�hZ8X��)�z�����"��e������+՞-�.������m���zJ&�~�;��jl���`��JyEb���gdg�
���PP��s(��`1+Df�z�D�0���2}y~GY%�?[dH���y�fGã��ũ�j��N��\]��"��m�9b��@�#�G��ɉ�`��u�4�x���ȥ����otj}��+`����P�o�7�5r�G:_Q��Uu�Ёh�X��e�`�C@i{��x���r��8��N�l��Wc��G�h�s/#����
�^Y"$��M� Y^�ke�v��h`j�����H��$���8C�,��]���g���%�uY�|:m3øs��3�d`E9��tln��T���lC�jB���]��,�6���Kb�+�5e������˽xg�o�%D{���f�R|��Wus���U��x�*}s��SC��4�P�\e�c�>K�'�js�����$�U�ϴ���!�����>*�٘z��}hp�@l�Py�a`fƓ�l!�_��9pt=*�u���Ԍ����q������R��+�4_S�ѱj�����vZ�J�����≼��G63I��^%�tFgb��{��y�<V�����V�]������g�>�r�5��M�G��!��jl|C�!V7I�dg>Ӂ{�#k�״��;T!s��(�t���ei�J���Cw?��R����փ��;���D�f���]l�C��6������,��~ﰡ���lp�؅^c��sB]�3�O�ɥGP�I�*χa�k�����S�p�!/m�����U��O@�N�a��Ff�w�9+���gv^vWs:�u
n��h�6�!s_#O�~E���t�Z���Z�0�狉액#(\�n(*Amd�FJ�pvX�Y")Ϫ>۝/W��U��p9$$����=���81'�,y�#8B�:"I'!:�|>&�P�t4��k�H����[#A�^[`C��@�pÚ�����h/(����l�W��Ǫ�j"t�0$��)���ߒFx�m�)I1̩Ј���;�y�h35�D��������9 ��:����>�F-���S�Q��a+��|���u�z5��Ń�v;�q���ٵ\~�*F�;�.S|̑Q8���DN�D�N2
��
msX[i<��1@�B���
��A�2�髋I��J�1{�Ҥ�ܒ�<ɨc6*�i��#̠���(9���>�+���\�y��`�]���\���CǑ�)v�jW)z.���qb�yFa�rak�8�K%{"�u��զ����I�'�����a-�m�^�U�ɣ6�Y�'��9�CLċ��r��B����uY;�/���+�0����
?@01��v2Č`@�z돶�:9��d���N�����a�5%sg�QK-W+̷�1�[�54�;j*d�ױ��a�N�c�O���\�s��Ʒ�ů���u��zB�g9}��
`�BOv+�W!�2�e�n-Cط����Y*�Rٰ`,0݋*�v�ʙ��0��5�*O����W�����������_��fye�)�Y�	��D�o�C��*�[ ��V���Zt�oL�2e��8�3�~�5�1*)���'�j�0UKMظn����L���/���bÂI�R c�mYz��p�w��>w�����w���� u��p[� �Թ	:����tR���v���1�0
�b'���(���q�nn�&�榽c8�@�Kϒ��ɕ�����=:O(0�7�#P�h�I�SQ��R�f�6���s��W�!�s��ބB/L��u��u�nG<�h�s�a��Az�����W��ߛyp�9�gvt�6���[ڔ-`����{��G$i�����e��6Xy��ѣ��PMj��%aʾ �)J���#��ֆ��w�KDq�0!�F~Q1�Bv�"��@Z��O$4�6
[Sf�A����U-�fk�rW���*�X6�D��<��1&:�}0T�j�v��O�P3�fM+1�����obO���ܶ"��ݢ<�o���A ����G5�Rs���KG�',�l~G���|� �Ѩ�Zb
l�њL�&$����&��.�Q:/�ĺ���g�`
h�[����̔U�PRe ���}�h�Nei�g郉��:#̅LY�*ׅ�_L� �S���q�� �ߣeM�8<a�.�6� -F6�koP����;�	�]�^C#"b�k�d�X�NgB�⤐��r9z�}���O����>ǵx8���ׅ9��w�G.p�_�U�"��;��m�(�!�m��o�Bj�������AϨ�J$ 8�~��:jd����RE��6VE��ys��[s�N֏ �1���a�-.�+G1L����z䤡9D����+ɅI�~�xf��и�.��2�[���x�yS�}>p�����z�(���e�+��Ms�80n�b��C�{ʜ.-a�onPUEB�$ۃz'���� ̎U���j�T�yuv��P��e<��!E��dŧV�/(��,zQ:���$Z:�����TE��ρ���b����zݲmq�w+9d b4�������cb�P�)��.�c|z�ͦpU��@Imք�I����&L�dY6��`c�M�/%	�����d?��v
�|�`.��XH�T�	b�Z���7�y
A�A����%V�9]v�RfK�˕DF q��*D��+�ُa�̚�/����n���:<�ĭ�����>�� >3$&f�N������4��U�#�(O_�8�q�EVR��A�S4��=�J j\���	$��t��l7�Yə�nBm�Σ�HN�j<P� �Z&���u���:�1Aʔ���,@����*5��|/��Q�]88��q b���h��_,m�y馶��=��z��໧3��?����B�hcPB�\�4��t3g�$�������p�ŗ	�5Xŀ���%Z���4���i����I(C�@-�2��AX��R�V���B߹{C/��7绲���0�4fa�+ӑ��H��"��l��`	zL0��4#|YY��N�X�y��D�>��
�q$�/�¡W�:C�@�e�4
7������̠��,�o�MAN�����|(��~�p@z;+[y�J[�yN�h<(^�q1��`�H~�0�������u,CN/��K_�,�� �*>n:�}�>n�l���7	��_��s��'lNL��Y�g{F��4��DT��̼��&+����o	�hfZY� �BcSl�ʾ4�0}PO�F�}jQ��L�{�<��W�/�vG�� X����yi�`f�2@n�qK%Ry�:�q5�|�3S��rN�gc������R�qv��Ȯ?��{��j�E���U�+q�(�9-�<?8���V΂��*�~;*�K6���E�x8��[�>J�C�M�\ɰ�ni5����u�N��Bhp&�.a���uiJS��`��;��x����+TV>&�G�q��{�Q>��i]��ɿ���$֐yo���'n�f�פ�n@3�"�d���b�a�S��6<�k��l��1����=$⳹Ly��Ŗu	����q$6��f�.
8*6���u�M�u�*]>5U��.�����k�����U}}�w5�­D�H[�._��2�T�K�`�t4o3�
Q�dK�{X"��d
8D��r��6	��eߕNMm�ہZ!��; �],U) �ؠ���{h&a�@�d�M��j�!񦁪���zfC4�Sk�A� 4{a<g��OW�ߘb���7>��+�E���z-2I�;��2�Hw�������ѳ?.N�!�I͚+7N�@D�vɖp��3�2����I��}��qa�S pK�`�%"%�3+��6$[���� ����V�y�����=MY�|34�s��]Ļi��@���pku�rwS*+�?�E+��V��&�n�x���F�+[*ł?X�+�w�ɒ�l����ˊ�m�i����+pKZ�����s��,
�H�
�4�L��PyL���im���h-]$��R@Y��J����_#���_� ��ӱ�7� �h�Q�T,78;!F��p�΀�!����L	.G�xLd�<��p�YY��D����!B��n2ҡV�y��_MaG��vń_1ة/[�$֔x��{�#�Il�� �J���vEI��J�� `�0��q�G˧Hj��TL�ʝ�ܫ@������k㖽!9{��ۑ���6��}���!hd�h�\D��b&����#�
~0E-q���x�Tt1NiI����<Xa`B襝l�����O�=�	�v���Y�rҜ��wf��F����yĺc�eFĈ�G>ќtx����
��ʅ����y����-~���emlۑ�w�&�z��6|�>�'���S��~!�	���	��%�x�w�&�+�h(�T3�tkY{пnP��\����G��gz�gQ�6'	W����U�{�*�1H��۳����Y���E�5���P�oc�Ң h�g�ks[�����3}��PW��ZU�D|�������X8�����]~ՠ����Ð��kY�3(��\��*��srj��d#/R�!��J�ZE	�".�Wo6魻#���X%2ܬm5ߣ�&*	��(�
���J�ٍ���lYf�=y�݆s�强I���-66�w���2,d+��~�E֩"{��d0����H�¦>o�e�G8���.���GR��7���TJ7 \�����!cZ/ �3���N/�fg�6c��4���B;���SF^O]7W�Otr�a���:{�\^�n=f8l>r�UB��94��Ε�5�#�qLZwF��h�]�]X��谹|`*�^jd0x���,���#��vaTꑪJ���{�4�Hu��Ȭ�-؞)5�DC���>T���Q;�e�M��A�l|+w�^�@Zs���ƚ��Ph��p~h��˓a������"���N�W_���"�U��d�[攐?(���+zO���oa��w�%B�M5,$�^��{n�7��f�`p/��N
�Vl�_�q�����ヱ5P5-�rX$�':%AOB�o2�\����c�Fu�O�Y�B_��
W�ڔT���co�c�6��?�����,Z��r׿�}�>/�U���RR��)�M��;^�)ѬE���?n����%b��u�-'� �<�R?������cm�<��{p���]
��)����+�u�Q��@����J��/�.��\�&���	�+~c�g�y��ڌ��5G��q)�A���b��R�o�nH�to�*��zU�Q�wޒ������dm6���y*��:<�̔��X���l)'�Ț�C���Hf]GPy�R׹�넁Mf`Y��m#i�֏��$�-��K��j)ɂ���Y���#u�%��1s /r�F����\U��~��ܠfm7���mO�K��O��ZnZEH�0{1u��:+c��Ah^�	!?�y�ӡn����������z9���}��u_�q��)�|���"�b�=Gly�J2��cm���������;�g�~V�.�ywd�_a��pSK�H���ah����U|�z{sjO�1־-���'xvo��L:�Y�F�+�2�P�ڲ q���|f�q��55�済ܩ7������F��;h����L<�'�P�)�*�6j�R�h1	���}��.���rfG�!l¾0ã����H;��m��EŞ�OT�Yj}>��}�
��!���O�w�I�JLr�؛4yV������6eT�X��j���F��I\�>��p�T_T��y��d��qb��w�6���7G��
%�yu��?ٳ+C�`LшL�5@u�J�f���_v�n���,�e$\�x��l��?\��MA�Үc(V�jʶ#7C��#*h�8��1�u˖~ajt��GCԖ5�p�F�8���/6[��2������'�[F���h�tJ�X��̞%�dN�i��[&·��	�?�2#��$h��V,�蘗h�h/�7_W���v��R�n��R��K$2�]�D�r�a�ߞ;_�i�s�C|Gs���� PJ� +�0�h齔�75w)���O�,5"�39�
���}�lZ��������Rۨ�ɓ=Yٛ^~����z5��گ7p��W�H.͉a�HG�lh�:��jȾNQ���N���y���CЖϷFt�R �YSW<����;�F��.��cMU���`_HgE�XٖS-�ю��8,�f��u�u&[d�@C�zvZ��Ϩ�!shg5�B������U/�����������w��C�ED����P�<��Kq�AE^$AuTLUƻ<gF灖�m�
��f��
	�|��0�Z�24׽���G0!�:�@Y���]�9�8�`�˾U�͈�,R0�'l��V3'ѬAr'�D��]��K��Lѱ
�`؆ Z���GX�r�Yj(7�<>�Y�)_hF0���x�g`+k�����%��W�[E]���F�@��/�O����XSy�8����j�[�@d?r���R��n~�;���
�%��[�Eb&��X�"g��פ��K�-_% �b��E�b`X;���&fN��� ʏ(�y��FQ�
����6L<�����zz{~I�4Ę����)�#k[!E�!�i'��F���a"»�$|��	��΀໋�ۧݝ�1�bT���l䋯���%���3V��:�[������|��G/JP�X���1���T��
�.;�-�E�p�d�	�j��6s'���M���*�/�'4BY�!t���<��'�Q6��Ė(V
�0��:�,��V��,������Y0��x�cM��#q��ӻ��(�U*�I�8�LRbi�"��S��o��}�]�|�U�����\Y�f�}U���o+=D8�7���z� &��W�P/��u� �uRo��]��e1��Kw@���CРv�X�丼��MuغBk���7� 0!j���?5c�o�O�o���,=h&�F=m�k���|R��f]��+�x�o�l�l����o����tBJ�I�M2�G	pX��+�Ǌ^s`hB�@�n�\�H_�H+�E�+o��.�ɱ���N�u[#�:�x�.�����򦦬��w�v�0��0�^VR�e�ۑ#ۇ�֫~����Zφ\�нU'l�l��@���\)��C�}?�p�����vZ�(gm*I >7�|݃3<vHB}�ϟ�Do"�{����O~�̎Æ�.��i�`/����畈�ԧ[���|�	'��:�ڰ,�"d�P���J���$-GD~�Н����g����u2�k��x�x��M�`;�����/D�O��֩�:�^%�ô���ȑa�:�ʦe�rD-|�P�7M��z���E������F� ��<�灎@gE
���:�x�D��>(n�s$Rǩb��\�S�8�FԈ�m�M ]`ǃ�yW ��]�d��s�D�)�+B#`A����f�,70���k��߅��A�e��7�B��"t�d�$��Q�NH	0i=�u$��vtjU�}W\��A�<�)��Fɺ�@	:�n�9�aN3T�}��Jmv��#K���S�A0tV�J\�8�OD�C}�$z0����l2I2��Xm����+'� &��F�{X$�j�R��O�"�X�0�����	�>.�,d����-�Dg�4T�Gü@精�u9�C�W��w{�C�{�\F�r�
�`�Qi`l��ǲW�����t��O�(F��^�eށ&��PF��Ƹ�
�&=֕<�Y��sa���X�|�bWFf�s�x�xs�%|�ӳ��W����%r��d�Ҙ��P\*6�����t:�~>�� e������k�} NЏ1�"[G�2�gX����ʧ�30o|cf�շ��
�5C� $�2Rz�Y9M�_� =�0K�zS�Nj�����2\�U��������[�SͨM{�u��/�X��5������"t+�sq���n��S�.��H]��Y/���U��A�X
/�����M����URof^W�Cx{
�4���';<֦��H��]����銨�7�d����\��d���ڦϿ�����C(�X�
^	�F���Xi v�yh(pչUsG��N_؞�9���h����j�2�Ǳ�L���79xG��9���#@�ɽ��$S�]m �A'�|��Vr
=Y���f�O`ǻ�ƒ>Νi賲XB�� ]�{���l-���'�A�� ���ߗ��/�;�R!L��q�&��I� ę��Bm�;�R"�D�(,�������p������f�k,�j>��ǧYf�w�NA���5�1��V��]0���B��{�x!haFSY�d��.�T".�V�b�\�s���-����;Ap0u�IQ����<=5iG�K�_^S�vҭ����&�{樌J��X?��s�}f���G X��}ְ�<�T�~%t��b3��}]�@�Ϸ����з����C��-R�q
=��~v��<ReP��q8���Pձ�(Γi	���+�z�f�;��"��8T*3��7ȩ��Y����0�K�$^�$!���o&��={H��3ң`���5��u��
h<�o?��|V:!�I��=�X��1�!t������� �⅃zV$;BB�9����V-[����J��(��YB�q�(�0�o!͟Cr)�<���t��G@>��T�%���%�n��ずz�kD��R��v<P��石K��^�	� .3 �T���m_e8u_��c�c��X�v�.�~[����L\��a�ԇ��l�$jx d���o����%-���Ɲ���>�}A���	��9�=�-qe/�N:�B/��)C��)(�`��]t\JYK���V�41��	J�%�,5;C9�J�B�5��O#
�v3�}�r��r�D&��@r��AL��+Bk���`V�#a�@m��0|B�����(ROPߤ��X$�A�R!���(Ռ����󊼨6*�`=7�����7��0;VF���f@	2�`g~睗��Zb�����G���N��D���$�wnE@�*�n4�(?�}������PC�HB��LB�ŉ�w�q������m��	⾳E�J��=�m1
B�u���lp݇e��@�Q_O�r��e;�$Qƺά�5�H��X;�����O��.�z�n��M�8��A�_�U�9�]���6�/N�v�a�CEU!}���#�o�e�ٟ]ƱMd�p���֑jLD-�,]���ؾ�	L�j� ��	D�#Zx�TR&LP%�.Ɏ��؁3���y7z�f���
,�W�?lH��n1��;p�%�p!��ā}/��a��n��̽�Ԏ|Ӧ�?�����q�w�K����`����;��cpHN���|���I�
�}U^<bon�+�>�r��l�7��3�ڝ�o�|:�.�������_�Z)5k*��2@e_L�H)F�nc���Y�����Br��w�5����>�`0��͡r���j1C[�l|� ;,C�@�
�6h��<"���x���>�!v�β��:������e�);��tE�/IJ�̗��J�<��͚������a�1h���t��Qپ�)���"��-$ø��aWw��Qzfu�$~�t~��Z��E��6P�%�a���uT��l&�h��mo�c���b�p_�?�w�}NE�i�510�Vr�N�Fݯ����S������6�C�I{��Ƀ�7nk_����bº�Fm;n�˸�QsZ���}����&�47w&=ݘ�<�|�������KN�X�:�}���T5�U
`��T	�	�ΰ-��?��8�ims֛=��z���l����sl"���X�f�,�����z�+[��t��/h:�x�Q��|��HW_�É��e6�5��:���H��I?� �Y��S�7 j��)2�r��h�;6Z��^�i~H�� �i���n�Ϛ%~ N-�]������V,rJ`a��R��[g��0S2�ִHa�YݯK��
4zB9r$�j��#��TpI���n��@Ϸ�o7X�6��SH�Xء��. ��"+qt��ӭ3�����=i��L��y��g)���T �j`Qt���d�K��+��^��d)�4�7����Jqłh�Q!�K%a�`�2����!��wX(�{Zۺޖ?��7�K���k�Qֱ����cEm�5v�x�{ITȾXfq#`��!�F���w
�a�@x	����/�r3�� @o����!zx
�':�1C�
zS�v�$����FU%[�m��w욵$<M�p���_�G^qN� [V�ؕv�efMX\���]�X�-�D�P�n֥R�:2���.��I���71M���(0��c<A��i��g�!��"���ua\��Z�����$+˧G@���za�9Gd��k���#��_ �8��z��ޭ�I�L�����[���_ -���4�ۘ�{*���x��Ȭ.����U�zl���^m������#�e�"��k7�W`��S=A$b�_�,&��P���ɬE������ys��΍�w�}wA���v�t2�^�Yϗ��/�U�v���ee�����kㅬ
��\̀a�9���r	�;]h�'e��iB��|����������EF�^޷�Sw�Ō���p%n���-�o���7��Ua̹��\~��pƢ��t9�YP٭�r��,"����z	��Ef6�5d���"ܷ"�;R��gD8�nai//�	AN��	u��F�]m��9������np�TL*��&��0�Mk&A�B��n]�K-v|M�'k�"�E�k��k�+�g���2��r�`������0�R�< �aP��;�o���ض׾�� �?N�{����$� ������U�+C���[�KzqMb稬"c*�/�̏�BIXCg��:��üF��EO�|IM��-�|k`0.9�����Cǆ2Uq���N��JHa�(6x	JS�U��X��G~b(��
Ē^� ��K���/�F��>��U�J؀�G��ƛ�Dú�|,tg��3��^�`��R�(s�B���"HO'-xw��x�lLj��4"��*��`�H"��`���>�;�ɜ Ŕb��d�k�d�5m���U<����~)r�`�i��\�iW4c�pnvSa�A�:��J�@*rڿ�ȹN�L�~g��K'߬�{��j��.J�zx`�L�����N�֞d^����ž�)��^�(0�E[7;�_��T1g��n���ܠ���>(��{{\�^���T�=nO���ĉ�n�g�.aմ;��5T��kx��W9�8A�/�X� D�t:zM�yp�\Pw����@\qLvF�ʤAI�ڃ#���&$M��:FiuI����"�u�.�4"_��1P[�����,H���ʄ}��5l>93�kji�e��V��S
^>�qQ^�4�p�ri��z'&Ϸ�g��F��M��v��A�Z��%�8)|?��N�2!n�MX��' s��\6p�<��J�*ბ���~�O�kx"�Z�@ ��\3���07�&����}�� ���|� =f���
��]ý�?W���⮒�6�\�Ϙ�(�B���q�W��0E@_?�j��������W�x�T�:�ᘋ��r��V��"�EQ�9uK
�6�B����u��L)ݗ�{y��.W�R����{L]p�#C��Ã8�r��E��N�soi�Q-j�U�^�~�J/�c�AĿ�m�K�>��[=1�� 1Sɠ���Eq,� �2��Rh�V����`aai/��S�#��^-ek��Ǉ�R��Ҫr�P��O�b�2XY���g�mZ�����h,)\TU�{��e?L�x��O�sA*�;�+��-��=kv=bi��@��&5�S�+[Kv4�*f�\0�>ѭ��\�]�f��5yh�������7Ǒ�y���CvPĖA�VZ`�u@�>��wkt�wI0�k
��,��^�Ӽz�em��U\o
B��Ӂ���� U��<�]xW�
�������Gbhσ�xF����M$���$[p-�ؖ]��ͫ
'�`��W�Ӱ�d����s�+���c���a��Km�{n!z�%��9����S-�ޕ�s�ua{D`���i^h����?<��	��K"i�Rd�Fzft��*��GD�Mk�8�VU.�bmf���v񙨱�0��sÍS�h����Mv�A]eG}�{�+8�
w���E�b�[j��jjb�SO�Ϋf�'?�4v�fek�� �d��ߛ*��
�������� �ɟ���\�Y��������=-�!��{K3V7�h�G,�3��,zn��2�����UJ��/b�-�c(�Բ��2�GJ^�y�W������6�$��E1ÿ<�Ie���Z+�3�f+�g9FHJT�q��x��sBĈZ����,<;��̘��Z�H7��`���n��mCQv��,[�#��D��,u�i)�ȥ�6=3�
tY3s܄V��Xb^�úշ�|�Z)�y't�U*?����B@���3��Ky��±U��g�,�}��t	�ŜV��3ܻIZ�s(��nu�^v{+Q�`gihC�r�?�>9�u2�#�gi?�H\�V*wG޲2�q�	�ֈ&�]<���JȻ���3Y�C��:���]t��*%a/:e�l�t �	��]kn"d%r���L�~�c!vIWWx��L�nS+-$1T~/*&�V+J��}8����F�I?�w*-?]� �4������q5��]�_�$�5g	�ɓ��>(\�>3�;��Te��#�(�' j��7K��%E]�<'�l�"^�Vg��yC���Ƞc�_p��a��Z
�c�H���i��!4G�����x��˭��4ƫ$`�
B7�c�z�{�N{BB> ܶ��h[71 ���������^��a�e"��{hws@���
�q�kQ0��D�)������`���5Yz�P"=wt�.oQ����/��� "��K:j��uz��V����>�b�oIB͝�S����
Q���������d������ݶ�)h<���=\�o8�mܗt�*���Ap�V}`�כ8,ֳr��I!�4r���GR1ֵ@M=3� & S�Lz���E؛ێ�m?��hc�����V ��~ĺ���Er���}�/$�fퟶ=�Uե�1rk�Ɋ�%�3u,���١��o�iU_�V��rS�z����z*Ct���{�;ڃ�Q��l����L�;�I0J�����(%.� ]f�d�P�C�:aL,�Ѱ�2[橦�BO��6�*ݘ [M��wc+�3 Q9)R��
�dom
����XP-�� =:�C�����c)s��
�<*��2�t���1D���_�����l�{H7D�L%��j	Z�Aw��-"��-�~A^]t���6KU_9�3�=bs���ߒ<�����j�S ���Q۾�F�?'���^��E&Z�r�]N�F������!��� �*ጾ���5Ck�gX�2����{�2�Y[��jn.����?���k�<�ņ�d�q�&�aD=0�H KFWѲ�7f��?�n�Z��%�NH����nv�	�W�v���F1d�p��뀲�`��. �;����L��Z����v�q�-�gy��ޝ�SH�V�D������6��[�����Z��Н�=X��P,�ǔ���	��4�0�T�ǳ�����]Bw�������H�|_<Jٍ�b�J/{�&�pҏF`�Q_��������g~��zD��;쯈U �����*�ܜɌt���<��*�ԲО����#�Ȫ�4����hi�V<�Q�嫂u���Gx�F�RU[x$���� ��O������/��h̘\)��a����+�{���2��^��ܞv���0u�GGd�,h����܀��xgT���F%.�#�&!�_c�[S@��^�����7�x/�b;A-@D�J<�qS��/�$�y�zQ(x�ntN0�}���K ���©���E�{$�.l�Zm��~�P�^z6|ʧf�}��;� �+�1Y����1I�߱y�7��e,�ARha��>{��Ƴ�i�"ÃR�V��O�1��v'��0cR�^e���+f��K�_!�G�����ph�5X��%|��`��y��74_����Ч��QY[cLV��W��uYY�F��!�;�Z���|"�Q㿕��l�Q�	V!�G6��Q:l0i/R)�+QҘj<��Gn�*����><���������e����<�#�O	���D�]��7x�i�����#��}�Lx;���ے�0�T�'HĐ�Y1�]뮌�����*�!�2f���&�%�}���4����g�JL3x@���4�=���Bx�e4\�
R���GL{�:f=KJZ�\���� �vư�!�l]��A
�W�ˆ�Ltݖt���c���
@��L����=%�y��R]��)����H���]��~����n~�0O�֌J��`�p�f\�^��ΰig���q�0c@�J����Sp�{�q�ŉ�i��ld~�+�(Nl�/��.��&a�VX)6�������>t��%m�o�|,,�@QI5Y�ufu�)�>p�F^�J2/0��t�~�L�n�U�{j�Q�@��ҟ�:�<��e\�~�0�Tp+l;��P��+�J��(f�a��J���m=����5�O�o��p�h�*Scf�S�`���Ӎ� �_>�Ñ�8ɒ����.�s��c��z��D����B�����M�����NU��*�#4��{Z/!�Y4?��0(,u�v+����\P�i5�K�.��Z��s�J���Zu�J����"���K	�2إ��J�i=U��kZw�{i�1D�a�Mb<�嵻
�̧��1ek����Џdpwd7I����9*�� ^������_*깚B�Rj:&�NJ3���_����)���G���X w�C�ܧ�z'0t��@�g�x"�����5lE���\_'�!���~Q�4)B��l�W��ry�'��>3f"����*���D���P3���v~t�2�`�8�'�R���"�� ��v���v(���Z,�:�q��T���	D�b��,����Q;m.D*��>Rڙ�Z�8��\"�\q��&B�*�F�|R���+}mnA���aUUR��)�q�{�s���l�����F����hP=@+ڞ�%w�-V�,���V�[���ۯ��m�����̜�`Z���98���_ǈ��X�:�E��uXq�B���s�2�Y.��ʐ.X���M�蜠���b���!v����M¨��7����]q=��a���zAc
!E�k��JZY��E��=�4�$�:��%z��W=�|��S\F�[HcO��nD� p��3s����Em쟍Oe����p_�S�Η��=���ϓO�6���CF+�+��y*3�p#?�P\�6�b�C�#8�_3w�m�� ���r&�쾥�L���J(Y����z���<�K�P�g>`\<��gI��ln��꟫����4b�Du�>Az����+�g��a�(��R��D������|V�F���si�u��A��5=�P���(G�B� ���f����ӏ������8�t>�{<�ڨN!�'NQ�Q�-;-������VZ,���=!���k��xL<����c�'�UT�-�=]J*�öa�v���3� �)�����::�j���ͷX��2mHW�=@�����[��TE��a*+���{]a�4G���N�o��ጝ�mO���?�.��|�`�@~�d��R���0g����ԥ Fs��O�X�����ә����}q��i"�����Z��v&9zW]�HR@:�M�͂���@��G[�� �<X��e7�c�̬�)<��(�.b9���od��?���J�R��S.4�-*`��0�z�K�`@�.��Q1���k�{e��8~�����ט����fB�6`	��Ưn>�Qo�,yf`4�[�G&���Լ�=ڀ�E(�CC�F�p�46IA��LiZ��P���Tsg��dlUF8/��M"�E<?��Zb�㪝-xj�k#���(p�ʹ?� ����k 9���+l�I��G�� ��Q��V�(�?ɽ���4��������/w�o����I�&6=`���_w�<'|@5cy�d.�*ѕN�@Y!ltw����� �-�ͯ9�cU�z0J�u�`�0#0e�l�Hs���	Aw�)�q�6+�H�q�h��&O f�����Jm��f�r���j;B��Ƴ���K"pvoz���"4k+p�hbۜ~���JR���ᙟ��@���W�A����Ba��yؓ����%Q]��u{^�o����V`Zc���TS�.}��]�������OLS h�9��ab_�آ;�R̡�w$���?�n�����~,��<��͔�{�E��F���a���l���ESY��Р��X��F���W����+av9E>�7�	�o5��o�u�a)ݦ:~\��<vI,���TѱQ�x<��xE�O�{ˡ��C5:� x���ލ8��]�\���OB�u�|�����|_T�@	tn�>�p�?Q*Y�\�_��hǊo��C� Bn?�v
p�)���De1u�{�y��ex_���Ph/T�R^KS��0j
�������<�C�o�8����|q8���}BҞ�(�p$�p�]��,����&�o# ���frh�ѽ�yBQ�⼻$��Ke��͕:;��������σ���������E��C�0��#汻�C;y��1��t`x_z䞴��P��2��)y��B����gY1>`s��� ���a��|V1*V��f���Oh���
U���q�c�
:�J;��z6,`����g�^'�&p�&z>��]����,��^��еm:���cr�^�o�
��zĖi�=ORGJE2��j��6����F���͒5��%N��1��b!��s�6:اyNiGy;];��j����N�y�qݻ��F�<;�t�U�Mh>!���W5]�a�r�$v��S}��(���������~�{�ۍA���`��\B�-����y=m�� �i7����!E��������
	���o�n #�>L��e��zC}�F���^D�p#,P��d�M��c@#��Z� �E�ހ���m���GI�SGB ڬ��'�٬_�s<��]M:.ll�{��?��?�E�����{�|W��8]�eg����c�8:v�������j���҈*�#q�'>fo$���y�hA�TP5�7�����pô�����qE���,�-f�3�Zi@Q~��~��P�㞝��~DYJ?:G�P���y����J�j�a�k3P}�����d�<s��z+јK���Hs	��� �e$��m�z��2���t���;���{#6���k2E�Me��Y����Ed^1��8_�;g���&�&�oh�Q9ߕ32�=�^5xn�����<>U~f�n�P�bU�נd#c�J��xPo���-HdY�e��L�k���f��F��m���]\�>���W�����5�|�a�+�Jnoq{�kI~�J�%Xꪦ�1�nQ~<�F���}�_�ܬ����D�A���^�1���aⱁ�=����1�n��5
�W��Y �-s
3��>TI-�E�Q+<��o-�~s�-�{bY��}q1�a�m�hLÇ+!	���2����n4?,[�9�I�-��U��W,�)� �'����$��g34<��	1~O�����z	>�^PϷ��z0@�+<����+r�S=����B��+BС��AM��5P��R�dj�ĩ���<���:��ְ'n�t��M����1h��.�
~��0 �P��m��I`	��ꗖ��$�7��\Rx�����"��lX�J����+n��=pp��/�Sc��������¬]�IZX��.�G� �^�;*�d2�Ո7M�����K|�o�v�����,�x�]?5��_�kY��;�+E�&h�G�3���� �$�F,	��K��4�� ���U0wI���[S�	�UbA�S���γl��n�F��8�ܯ(����Ĭ��q{���N�Fa=��+=!�|�j�O~W��������Z��(rܴ�9o �/������,��A֡�S@���l+�vv�t��������] �����1Z�I��d�E��jr����"��PS?�#�Ь�=�>� E�F�?k׉I����1��NC�8�����8��J�O��>g�3���΀���dN����>'�6Y�x��?���~���\0	�n-�d�W� ZӴ+�� �p�@F�o��ּϽJΥ���!�ռ�O��=x,���$9�l[����1|i�k��X�ޮ����Wx�}+����D�>�� 05Mʜ�/N%ѻӋ7��ʶ7���Z{���.����!�j�S�b"B��ZU{x�����zx�Hd_���f:k����_�/�gE�-KAC`��E=���S�����0z���ufG_��ND��V�X�k�7�g[��޿Z��x�й'�����ׯ�ԬZ�d�?����dh\S�gu�/ ��E]�H�Yw�j���;�5K*�XBK�V�g��h5�B��)<#��fT�{k`N:)�z�X]�����.�-8�+v�_�8�:*�) ���@� p��xZ@P���9�9��h�@Ӫ�xPv��+�׶L\��i�y����;�W]L�m���ƛ�� 0�����|��M����Ⓦ�_!��/<����'��bf��{滥Z3*ww^v�"�M'�H@����I��mB�ֻ���h��I�Z.�]��$��$�w��*m��'��j�9D�����n��${wt�@�~�--Z��d>|�r�<_����s��7�d�i���e�1�t��֯�I��󃧑*$�7�Eza3��Ҥ>�9�E
"<��ɏgE!>����cRD��v��(u}_K����A�9����kn`�`��wFew6�j|1v]vfjĎ�N�\�H=�Ţ���,��h֏&RY�A<��𰩑@@#����������x�f����)x_�w&�fJs� }�_K(�]L��b�l%��Q?�����/crri��J��G���)*�_g�;7�	�$K1��L�O�a��1�I{��){�X��
��k	����3����9���ݿ�3i�nYϧW�\p��O�G9�y�j��+d��%x�͓�>��MӜa 󅏼��Iqņ���l�!�/�.��-�%�˻|J!R&J�[@r��|.������K��֠�Z[�j��A7�N�%�@�����ec���{k��R�IA�X,7�U}���b���.�~�_U�hI�b�����|�<~u�� 5��^Z&P���%52�@��0��� �n�W��k�=n�*����%�O�\��AU��D��KcB
�+������2��c#՛DL��4���(�Y��&f���d���\��:A!�ST���3�EvCe� pW�Z�}�#ݦ ��@X��"9ߞx�´Ϸ�]�˯M�G�����T��u̨"� 8͐Ȣ�l8W
8p�Kc5(���AI�j@o�*�$�������� +VW��z���\%	���bjσ	j��Т����}���Y�{|�t*1|]c#��Nd	�nc7���C��`�6ad6���Ñ�W����P�*�e(�8BF����ԌGc�ßa�`矮y��Eh��Jxy2�!s'd��֨�#1�����	�s�¡Q�gU�����ݺ�=�Iv��nL&�S`�ʪ� �[����vN�ܟ��$u=<)f�*ָVM��
�+Ҥ,���DO�>��������I��b�02;1e3�Y"%��J���u�Rb�zFt��w�`�;��0(�fg���yz��:z��u���扷.�h��j�B=
�)�O��!��!h���aߦseʼ��Cz�L��2єBj�`�� �=~xl��љ�Xf�F�EiU9KJ��#W��4��>1��@#.Y���}���uVh�卒�TȴΦq��l��T���W3+�+��'��q �0z�M6ƅ�h��!B$#X)���~>{���+OH;�p5J��h*��X�v�����<!}������po���i���/!���N�1��'���oQ��f�J��V]���7��̔���S-�v[���L�Q̖�TK�#I�YR7w�Ya$���畢����@!�|?���䘆\*�,��&/>��)���ƚ��4$�~��	G�n�7�=U�"���JRI�}K�Z�s�����'�k�D[h��j�M���(��j^��k�I{�M܂�5��!
��ן[+E�{��hJ�HS�ە"I=�����Vn�`�a�Q�U c��^�P!�y�{l�?�K}B/�M�=��>�)�u����>����i8~�a*R�hf���Ö�Z��Wｯa?N�j�����Q3nx֣D�a�7�S>m��_w��K�xR��`�?u ��J'o)O|71��"j�-�W�3����+H[��/+(b�M%E?�|�A���G�Ȣ��8���W(V{%��c��rpIܝ�u�Ple_��8$�F��<��x͛Թ�yC�Kᒭq�G_��DZI2����Gg�JH�=A�W%:D ���@�iAW,:�q0�����ҟ
�~�ܳ���� �I�N��9��WE�}���e]�E�V^w�\��C����0*�K�uϖ��v�s* 0�R*�o"��4��u�$���mD=�� ���ּP�S�3�
W|�x�r��h�Vl��(�l.4q�ˡ�x���lHoj�TSp�ˢ��jK����@"(�^m�!G���sl-�-Kh����LZxn�^`�E�Xq4n�*�U CX�ԝNڌ�>���3�G9�X�
q���W�&��/�O5�G��d���4�!�(ӈ�RL�/���pl��M�b�o%�ǃ�w�C3�����%_��YI���=d1��-$�j0��vr������@E��B��X�	�����O�yhQ�s"�"�G�e;ɨ�F!H��!?$�d�;\�`U���[bUǩQ� �s��5��4�SE�m�Q��1H��7��lRki��:� C��T0���R9zM��&�I�_�eV��ה�)�z�ϵ���[�J=����QU1|P����΄G�5�$l��#z%^��mp���'��
�fwma��f�>R��ɏ��Hc�wGϜ�J����B���IE�3 g�R{p�y�Z8��	K�Nxm�>5)s0�(��R�;�x+���Xh�� �Ӿ=w��0��={��BDVѫ���C�I�6�Ww>Đ�hx���je�������H�Q�V������@��h���{�+m9�V-��
HQ�ٗ��N�,�-w�����מ�-9	�����tv4��Nt?��͚r����(>���Jh'7z�H��$����?3������5�Z7�qF;9���8gE.;�>S�س#tW7J	9��9&�k/���4�� eɍ���-�)�P���.""��/����/ċ|�{(�Ip�Fc=��,�[o)��2�i�9�@��1���!Eg*�������U�w�J7�u� ~��'B��~2���#=(8
*���Y{�/�߅�,/i����.�	�,���D�A�"1iPtd9ʸ޼	�	��d��
*���*V����Z�ez�ؒ��(0�]���Lƌ����2�	D��N���(��D�j8��,YqĐ��}q:11�G� �5}-�f(V��?�;C��e[��k���3�҃�}mehv����1Ѡ��V0i
h��?b�TH��&�$����h ��&$^��f�8�LH;^�2���}�E`�����ɽ2M�E��� wTr����K�l��)>r�F1�UQ���!���__~���+%�*�a�n���-�wǙ���^�Z˧�)�b�9���	�\X����N�� fnSW���H�����-�WB5��f����-a2GX��b�\�{�9"5'����9*���^q,h�-��[9�$Yf�l|���#��;��4���ޑi���vmS�X���մ���:*,Y�	�N�ǡ@~�N9��/��.+s`'q��¹��!�Q���c
�|�dG� ׇ(��T���X��>�
����I�9��w�����3hs��#�D]�fp��5�r$�TP&o��2���]�*O�u������ui���vuаv�^��՝:M3%����Ixp�w�?���P=WI�\�Q��g���ᕴ!v�
�
Fv��� �'��p������7j��oD�"�Ol�@;�4)��K[IK�̥(#�>��q�x���G�BB���+���LH�S�%�/��;�j2�볙���E(�!5B��u����,d�-�[M�@B}u�C�D�� f�r�Al�T-9�s�eq����P��5k��]��u������т=���Ϫ)�|���s{�
֖g�bX�˟���	�ZT���Tµ��\��8��>C ���;ب��\�C��)��R칓���k����فƓ�țT�ed��M�����>���?ua���Wj�e{��c���m<Y�;�ho�u��K�į��W�n
�%�H�>�誝�(T�� 7�z:�׽UF�H�'����Ěrӿ�Gf*��](�KH�T�l��X�Z�u�^���xPVnH��f����$��S�WU�
�CC	��H�1��>5M���(,ё��r�2-?�ư5�m.�ձ���Wػ�r����p
�]�7�E����1L��5/�&B�0%:��� ��RR�!#å�e��e%D�Yan ( а~V<
V�����c���	+4�	{��������{*9?���zru͛��F0cY6m^��Yh���5��E��L,�uBPr�p�b{ޅ���nI�qO�U0�>K}�r��#E(�*�����su%�J�af ��.EƜv�V���@��-BRE�ߣ���pvu�Q��ャ�a'�<Ú��|G���E�S���d>������qJHh^ H�|�h�Z��zN�Y������x�PI���#_)�o�O�)� �Z/gC�W�j`a��N*#�X���#�����А�:�G�%�7�>�z���L��2ݥ>��ӳ5�YK�J�<�7���_��ީ̤2�s2�3�L �Ȼ������bG{����&�p��ŗ�ۈ�� �~���<
�vga�=��K�ݲ�-�(;�S�lc�����v�麦hCݲ�}�P$ښ.��y2Q���wp��Ӎ5��(�j>�u�|��8�C/�� @0����������zr(���NK�gb=�c�%%�o�d���n����p˚jw�i� 6!�Ɍ7�`�M�60��
��������Nm�>�o���]Uv�*v�)KK*Aj��gځ�D�������ʦiZ� 3�bI�����	E���;ˀd�hUj��A�MUv��a��fc$�i��Y�Ʒ���5�A��Njf�^���C8<#�Z�#Φ]^3�gd�Ŗ�!<�۾����Y.�!�[TA%��� J4O�����K�CeL��V�H4J�1�����;y��Cx�}%ꓫ����:�������a����P���:�W�{]��q^WyO�V�J�5L��I�y00����9��0C���txץ��b�:imԝ$�Q�~��Q�+�c����YR(EnGK����l���|���;S�9�Oh�;�]��tr���jE`�%[GB��Hbx���$�sxLQG3ҍ�in!�$y�!�G��P�+3��0쓓��t.�x1�ҿ�>X��2 �j�`��������X���B=�'��{�����'|�+饸���h�V*�w�\`�1	�%��)J����,�PYE}�@�S�6�.(�n�`�]O�0Z( D���杪8a��.SK��)��"	ʧ/��N�Oq0�3�{+n�uW��}q�D���(c��䪞«���
�8�_Hr����w�NKa���Ǖ0c�C#��j�e��J�yc�&���\)�%�~V̨�P�+5������#5T}D�x��/�9)��a��^A�gj`@���L����>a�*��Gaj�x]>U�H�-�|�s$"f��d��k��`n��+�����3+�m_��r�Ǭ�>w�ʔw��+M=t����t���� �L�a^7�#�ۤ=	H��E�U�^JT�.6�Y�ސFdp�ק�Z{f�i ����~}�XY{d�\\\j�Q�*�N3��Z�ϯ�p'�q��c��;5��![8N�-ǈ�.��c����h|M�&�'���d}tkM�< Lo��{eۘ-�w"��"����!��Ӫ>PuR�"zhdW�y�& �ٯ6-�撾������'��(�f6	t>8��($�#Aږ�"�$(`���#5 �x\�j�<���~b)�����$O��0�� �~����Fq�Ͳ�I�bH,���T��l�nBa�kb幙S&�軗�ݥ͸r�d��!���ҡ5��؃�B��"9l�.�8�5qR�7/�1b�z��xT4�f��{�O�,�sF�.s�IBx�b0��CA˫I�Y��r�$s?;: i�R��ݗ~Q���?ר�=��Y��mnX_��^R���]{:(uϻ�8OjMԨ%@� Zf��IӟF�\��t'[��yq1�';�u��w�Ԕ��vN����P�LU�����~�C���(���Nc+�0]5�.������TF,!�dal�̧���U�$��V�S�7@R��$g"4nNY�Ǧ�:�NI�	n���t_�E�ֹʣ~�fr�6�������s���b�Z%s�!U������/a�ұ*xY��\�G�>K��cn*˂����h��l8������<��/g�y#��J�d���Q86<�ո0s)�Y�DZ����Ȥ�ˤڍ��iP�S��"�K��3��E�1r���1Tʷ���aL�.G��� *�
��0��^��nL��XVA� �#�����b�����>���4���Mǚu°)Jx�P�F��'��PC�:و�����	8i<'9�z�Z��Vv���}�'��܂��SP^�qTv���Ǝ�v���y����P��a_�O��o�%)��#>&yݬ^�w����uӚ)��0���C����u�fK���2�@�K\�l6΃H}4�Jf)&)�:��.hV�]��*�0������>���U95����2�J�.q-(6�	�њ|q�Z:�%;6�S�/N�X[���m:�P�B�,�:i�R��@���J�룂5@��ڄ�<��ܘ��O#���EѨ���ȄU�@���@�m�P���TI�3�Ka�^.�ү����t�Lb�AB���`��>���I�P����
����d9\y5�hC�@�w�Q���M�~͠[���L2
+V�Xש.�	0~�Rm�;_�Κ#^8nmLE��D	F�<�2�c��4x�����o)����<P3	c�e��%3TP��6FL-�j�������7H��ԏGGv�8T� �QpL��K�2s٧�ؓi���;�I]��|�]�\��� :t�W���������,n�u1���7��
��!g*p|���Y�OQL��aÚ��9!v�ȶ��@����O:�f�[��7��:4�j���*�ݰI@�zZzN3�1����CaFmB�c���9
�t�Z

jكk.�DM՜��`�KծZ�z��Զ�h���Ed�[��5D�L�1�ˁ6��wi��M+�E<�g��Ǆe�=���W�72�q�B�0�n���	��_\=����Z�k�7K��8���r�{s�5_T�����?X4e�:~�"J���{�,�f��ܑ��ɸ��8�n��Z�=<��s�� �(�����3��`���	�rf_c�0D�N�sem46���!{PJ\��cN���
Upfa���Z�)�vZ`��a�Fӂ�Ң��ܞҺ��6�)���l�@�"gsDR ��y$Uxi �n�Paj!XJ�O���$2g�2�jc�*rώ�g���kf	V��"�җO(~�,�e/���XY�yu?�w?����J�ڕt�b�8�~H����d~Ψ��u�,��g�Ȑy���ٹlT�0u.�J�}S)��4=�J�M�	M蘑Р|�v����!�G�Be50�6s�p���Q+�4�^��,�g���
���EI���WTC��G��TC��=g[+Ib�=l�G-@��`v"�#�+�8��E]�S�i<X�0V}�$��=���n�	>���lCx}VU��p-ޮ��Xyu��w���>k�R��`��è��Q��H=K����X{ޗ��:�]���\BM.v��+�	l·�С���ug �1�J'W���B��X;�ly�S�3	������WT��(O9^ �����g����S���V����eE�=I���֕�'g�Ͷ�+�4�0���(&eYKI�$N��a�?]�{_�'U� �k�\���燝�Ⱥ([�l/���R�L��G�]7�o�۞4��U��Ƒt�<�tjllF.I������>&�-e
����xŲ���1��7y�c� �`��r|G��~�Wppw"��/8��^��?�����a+ ���'��`���,!e��u檵-ȔA1oK�4|�Q��;�u+B�^��
"��)`��D$��O�h���3XnQ����P�×��`&�hW>��lN@M��R�����1���,��ml� �,-N��.d
,�kP�>�y�lWyKh����7�4n��x�¾޵��d�cL"�5�U87hð�b�_�8n�_��xz�^L��y�A~A�������<O��ȗ����$��:'{{���9��zyDy&����D���_S����D��)ֈBI�.z�2�����J�]�����.����ן��2�C����a��S�(�pI�����n�96Dc�y���>d�&+w��Li�Td=���o����n휄q�E1�|�bu����begh�
�(�CRT7*�+:�:��z�sq�S�͝ŀ�uk;�~O*�Z���X�YJ�>�M���^I)l�DA?�UĦ��^\�dYY��#l�d'�z>�'�����X?y�COGk��u���U������5o�|L�PM$��}i5c��V:.٥NI&jO�%�y��y�4ڑ����C�SE�đ2����b����~��Q�i'zm����
#8ۤ��q��z����`�Y����A�1�xX"�U�)\�"��tE_AN��GFH]}��l��42�Ti�	VN7J;����d�I����	�m�Q�+�h�d�л9ym����+P3�DJ8tL�]�6��U��^,�����F�K{�4|(��#�JL�	~���TM�N]��EUD����?�+__{����(�o���Y����OR���cB��nx-��A8b� ��7$������6k<U`/32�j����l���~5Ye����<�G�^8}��[�*�t����)]h�+�w��)[���'װ \ܶ��2tq	s�&[�2�r
|�1��G���e%:j�C���̎4h@�k���7�FS����!�x�ڳ��_m�����SkR7�h��F�I��흇Z��nۓ�9t0��gv�v+�9�|龬���Ow��B����Y���ז���O���^#G~ݛ� �]��@<�X4'������3<�#�'� 1��[�g�T��U*�R�Q]�*� �O#�9�;�6/^ptZ�e�޵Gpe_!�tz�
߹���j�>ڷ��8�%΄z��!7[��f�c�74���[%�+��d;[8��p�p���G�� �Fl=���;Od�w�F�՗"��f+��[�*��0����E$d'��[�(��a�-�#ِnPG����L�,X�ž_��O�ڼ.`*���Ux��ϣ��e�Ac��γ�(�i�|g�ڟ��v���=w�%�[��`�[�m�""��͊�W�<;��������mǙ����nUj^t��K�"wZ���)��+T�-���(��j�_�a��w-<�2�XPks���#�t��>�1lo�R���r��Y�%i�a'YJ6�F�C2m8px��7�ς���^�����)c
d-�NI��.�/�c��X���x{�2S
�̑�j$:@��el��A���%�82}KI+?t��{�������clVY	X�H��E�Ŧ�[}_o���P�S��{ր��z�]��|���Ô��|J/9R�v sg٤(G&��ÿsq�c��[��`8��pG�n�=���,�'@��{qgÕ5�V��wE�K���XW>��1Ⱥ�I�������q�OO�Ԏ;�G�/
ZrR�t����TJ����'�G}�`�b��{�)��� �P���O�����k2�?[t{]o�t��jP4E�G��\E�y��
߻�Y���_.W���#��ي�����P���	Ub��
?h�L��S�v2�}�t���Á������X0������$ca�GT���ȍ�hc�����#�1{�
��]!MUDF|m�υ�G�ۖ�:cC��2ӡG7�.�H�U�L�;�9���]�5.K	�P�3p] �Ⱥ�w�a��٨�zl'2�O>�}�a랻���y�=n�B�f�-��w���U/�c�ES:4���?Aܺt�!�z�(IH^l�}������Ȏ�<�����?@�O�N7���F�ɷ���J�M�Ȅ�R��ec;��<Oy=�*.*��COm�1��p�<)��m�q�6���Vѷ1���K\6xf�e�?Vp�ӕ���N��#�u?瀁3^�s���́$���2z x���R�O��߷����/��+;K�B5��g�D��%x�ܰK�x�۩��s�g[u�j9�GY�iΟ�Z5�w���bt���5��:xO�J��{����l%{���eO��\b4�"E9���~#ufh!I��N?9�����P�948��{�c������:;�&0V'@ï���U���um"���62$c�V`щ뺆�SZ�<2+����B-c�A�L����`}�aw�M>A�N�����9zR��K̑֝ a�D�h��dp<�S�
�u �Ϫ����Л�g�U���M��q����n���R���:��s����L%-0=̷R[t����Ѻ%�R�j�TX��|0gزFV��6�ν�x��A��O����u�>�-pX�b��N�+5��M@-���xo�f��]��ݗˎ`��)�U���o��(	���-�CSsI��1s�/�/�k7��`�YZq�vOl�n���,~��ݙ�GA�3'/q�V�"�袋{epT̘�zMN���eJz<O;Ã]�4��`�o�[Y���m��&2�*�6��ks��S�]Ѷ3��F���_���"c� ��d=�?�w�@F�Xj�/ح�,m-��+rZP�yկ[%4`n��R+�@��C�b��N-ϻv�j��׺J�fQϑ9����}VklP��j��huҸ����C�)�������fh��;�7ɮ��T}�����e�D�bh��'�l\!JO�lh���@�a&��2Af,�Ao�N��S,<їGCEha��C���޷�����t���7�8Ф�����"�it�V���8�BIc6��}�e¶������LS�ZWh��W�E;�'):)(��R
%���C���11�&5W��u~.��f��M`�'��J��3�s׆�l�e{��k8_2m��*E~��gңˉ�{���]������H���4�%���HC�\;UߢF���j5sp�����+����$�Z]I[7��|���-���B&�d�Ei�
��ۃVZ�p�e�jD���{8AVoc�<&��v�att�~��!��&G����a�-��M�W��`���a�	��ۨBog�u�T��5��.���
�Y�vsⵘ����?�*�	���u���ͩ�N��O8� �&��G\�#��e
�1K�]� �*�	zb�p�%{M�>H�/�I�X!�H�����% ��!P�-��<\���Wn����=�i{:�@�C���I��E�D��LZ��'�b�������p��X荤y�R� ��Ħ0��X��*�K�G̄:��/��G<7ݱ({'e����O Ɯc8<6����W9D��u	���#%П������m)���3'������YA�?iF�"�s�澯��E80��춂+��:��N%@*�����<a�:�ȭ����3%�44�	�
�b�U]�̚�x��V�n�^.��x~�N�%�E��;p��8������%ޒ�����.~E%F�ә�~�隢�W����NS	�*t�pnl��1cbk����ɫe��L��n�P�'�f�dHSr�8f2�lw����e�ke5m;Y�M����\Qvp$r���#��g�^RFp����W��#��܍����3��#�=J7�47��	k�"�6�x�b���H������5od��CO%i[j�O=+��$)�TSY�Q��$�
���yf%5В*�w�?�MCnoO1�(��Tl��u�����j]()װW�hf��s��gߋ��y�����p�WZ���f�/�m;��,���l�@G��sN3,3`T���s����`�����Xz�h�>�<![T��W���&�����WdY��pIlrO	�p�ĎB�/C̻�[O�y=���A������=P�I9�C9��l"Wc�3���@�ދ�� tu��[Z�+k�@�W>)3�,Ͼ�0@�5_,��D������@�,�c}�����}gscr'7��-�/[gb��&O���j<P�k�ݢQ(��{��<CO��n�y�kxc_���8�`�g�k{^	�F�m�hZ\'�1���
ޥ¦�~�[�h֔���*�M����ӧPe��A��B��l�o4uN޶��v�������&x�z!}�@UOy�$�S���u�x�*���]�������#����|{��^2��N�U%��tɝ1?�Q���۹�-ߐ($�:��p�4�%�܎L�k(�F+��Z��0��nm[Ѻ 7��d��D��e1-�׀q��k�U9`s�t��(1��mpk�(s&����6m��UQ|�`����n�˵�?�[��M6�3.��JXBک��[Ěq�/1�xG�B,�o&�z��r�z)u�|�Y��5��6UNs�� I�li����K����nw��3~�����f����>�B��+���X�����b����I�9��~�(���h·�]gc�9���C�� ��՘qp#�7
�
g��?��G#z�Io���Q�LN�KN3�w�l�u=��P�㴲f=����#L�7��<뺄�'��𔶣@�a�����g6��ZK˩{�c����/�bB�����P_�J��s2��$J�eG�1�~̝Un'��6�,$���z�F���W��y����s�޲D���1���p��)�rm�׉7&l���-��N���a~R3�0�+��FF������C�?�ˊ��х�5��|�1/j��|�5��b"���I�Ύ�tv}�
ac3�"�T��WO���R1X����=u �v]^J�����,Ǘ�a��V��XyO[C���J��Sq�V�-�O0W���U�K���ڣ�)��Z��j���O=�c��H�a�A��Z�"�ޖD�((���� �*dc�",j�D�I"&���)�*:�ϝ�{'A��W�9�J��Nk�i��H:�J�ǖ���/s:xv��R�.��ZR�,�}���g��<h����IdZ)BTvĶ5��9kB��n���� @G�t(S5�%ι�1���9/o�y�-]���j��Sa��� ؘ��}�!+�v��޷k�j �<�'�!�:�~DcA�E,l�f��׫�i�&
hW��̃��t�Nl���ȓ���f�N������PM8&��R]F��i&�+~��^9O&iZɗ��U[eZ��
�����k��=8
Ɖ�T��zj8<�op̟�^ō�0��� �M�E��2��̌�>������L��k�K5´C���-���vU�rD�k�X����I�cg����(���˪V �8��kyN0�f_���������u�l��<���V3����;��=��x5�<z1���P�u�+f3H!���Jy�y��]�wBz�;q����@pM1ܹ�cp|'���孄a�nc��?�v�W���6��s��ɬ E���}�=�tREG�7��#��3�Z*�>ֆ�; 9�h��q�a
śXǜ��d����O_���}t��G��I�c�¨jk�� ��@8�"�L!]hL�sc�5Jl,,���Z�~x� �։�U�uNf�+w%�n���t�1��q�ϲ�鿟u�̍�}*�M�h�a���q��-��R�6� �z�>��C� ���#���d~��bf���N-�����+�,>4����X%\Gt��_�{(<E21�I����f�s�`����Lt(��#��k��'S��L�E����'�i_,���/,i^j� �,�����k�1*�̴�YB�>� � 4��cH��o�������C����S	j�H��������aԯ�����j*�ɰ�D��n�f6�$���h�F�g�r�����oq�����6ΈB����A缜x�]'���3w�ݷ�9ͣZR���D�4ߴ�;�r�r��e_b�-�),���e��8F���C�V/��JB��$P7
ZTt#W�MܟW᳗k�ϻ�->&�|���ן�����m���W|�î��K�ٞ
����0�v��ųY%ذ��8h[ܽ�_J��.�C-�����*��k<]9�{'=@�E�PРu&+X�_4+]Q(�ʆz��r�TC�*�0Ψ�`o�ܯ��\ک���k����(��c�J�k�Ą���ss�����}i&V�tS�;�k��/x���愣5��N]h|�{���x
��b���W��|ɮ?w6�Q�\?�x��[a�>8��Xr�&֌��x!Mz�	<�����YJw�ۙPs�A
G�*.�_�I8���smh���)�ٶ�UDE��cc�� � ��.~M��M��^Grw��b��?u^wzsO��a�+t�'wd�f�
�6�n�yG�u����i$ca�~f_��Sju�|�����)�W:9������/s0��$ ^�,�=��C�)I��^kc`P�C>��S!�1�.R���M�	�#.x���Ν%y��0�m�y��i|�hG���Mu=S6�rJ���uT���;��|₏�r���tQ�~�e�Ɲ#r�^�nU�'�ڇw��P�	dY4����2��=�|2��}�n��S,� �=�����7ע�8�-��hn'"����4��W2"ϨV:��{�g��F��9'X�O��(z��_����]C�4ُAV��ɑ�@�[R�5�tNy�JXT82׆��2!b9=��F!I`VK���(u�+`�A���J�H��O����lA�djR�w����Xr����H�:L���9M��ؐ{�
 C�R������J���W�f'��U��;$]a�����s�]�:.Ě�$rW� s2�ON�f��J�\u|�C���Q>{�kI��jS��;
�n(U����I!��)�9U��
t_J�+�IP�Y�w �gHZ��~μ�u�����a�~+����V�������[���!P��_�fx!������϶Ө�p��I�!���N�D��T�0}��'F�]�:_"���{���&!��)v�f���B���{e���7��>�T��^y�j�ņ2�l=V,z���^���Ԯ(�ٷi�?���t^��\��+v�W�鷳�z�TO�~Eפ����T_P��
����zg��S��iU��,die���mtR��]g
�F�FU�A����rE�!3��zx4Q2���2TU>"�&`�[�D���I�N��,��nN�-)"d{�y̞�;�WRDyA��c -�\'�u���)ʫ�ϥ(igt�t�k��ft\s�c�dZ}�r4gk�Yj�4!f��_�� gu�94"坛��D��2W��6*52j��>���[�| �k?"�Aj�q�o-V,�����A)��!��M�͊oKtҍ����j~��]�CCZ���z��_<O}p�3͡��?���r�H\ԇe\��b��S��Y��7^Q���x���L�"c���B��9���>� �
d�o|z��1���K>�{�ja��/��&�w�b �{؄�ߗ��J�1��P��ջ�����j��|J�"�i�;mH�!kN�0�a�~܃���]P*��g�w~��t^!dߖ�|#�ʨ����\��ʆOT*D���PY�s��6V#���9b�
�[��7�&㹎����,8Ꭰ���K�]R�5M�k�OV�	b��������3�<��~���OLә;B�n��T.�,d{����j��%�mؔ{������A3�ſ�������-�\�7%�B)oj0^֠3Au14�8A/.��5s�`��¡J�a���"ݶ�)���_�4�/ZEZ�ȩ7�V���H_u�t0HNR��p4�4���g�L��_A�p�&=�U��|T{�h>��$�Ȭ���$�g��b��BvYo�fh���a&\늖����M�<�,|�W�3���^��T�Xʕ3�_�ǿ���LJ����Ҥ�RT�%ǟ�I��N�Su��m��}Q�U~)PiO���ɠ�@�ܱJ6��2�� �A�7ɽ%��xK:gn��{[1}h�SSa��	��@��y�.Y)5CdX�$ѩ��^�Ϟ�տ����h���#��:o;qq�FT�j����,|2�@_)������"�f�	>B��}f�d�P sظ�͚t�}k&q�>���T���ya��T��2}	��2�fi�>�;���C~z�M_�t��?�>�!%�:m���t�`�F�2�j�'0��w���
���Q��KR%���2ZUƑ��o�s>�=Yu�%�M4&f�j__�RH��_�#�bމ4�Ԩ4��S�������4���#qn[�&��$�`�[(�~iC(�K�ݹ�u���s$sc�a@�>���&���F�Mt���p��D�Z Q����Tp#Y�쇃�pf�}F�C�S���`OR�(Q�֬B � @7�do�ߓ�G/�X��z()|ʔR��o>'�Y<X���˂(8��m�?��A�,���#�����u�
�2�
�u��uE �����\��Z<9�V(�"y�sZ� ��#-�+,�8_g]�m��F��[!FS��Q�v85�-���=���1�x�Z.��*��"=�p�f:`
do�j�C�dF��P��j3�p2�ǀ�ؑ��7\h��7�s��=+��	��8�ُ��Fu���/q9*]羂��&��#^�Y�A�5�I�{c!��;p���'�C��,���
%M�4�a�}uI�!IӮ��E���ڡ��c�2�L�dCmXo�|�>�4BZ(#��'A����0�JJk;�7Ӓ�`?���w�3����$�%
�@gQ[[��g���<X�d����[�J@TF5��*�G�����E
�O[�aqg$����
	�9�~���B��6,D4Wy���Np{�"�!���K���,�Xz����^������0�lB+Yd%�=D�y^
?@у�Q5&gA�;I<�Y*P�A8��.Q�w��Z�+�'�QF7~0F��V,L�b��^7R�tY��?{��YG]F�����|�9(�0�!ߡ|�B�Zll4?t\��J��6�X��<�Z��,�� ���8M�=G�� UQE� ����O	G;=TU'mM�>;dP�H)�TqV�G6�Y{�<��V���'ఋcu���[���������#���#{��� }�/�m���XZ�V7<k��</?�-v�Kkos9���<w�'�OOD^�L���4��cm⥿�<�Hx�^�򸹝�!�;^����*��	f�rzX|��^��;��L��W������ã|��=/y�-D����T�k�r�9 gYG�tE��jёE��5��q�' AR��B��p��ar��N׈J�K݅���)I��iJ��b(��˪�-A�Sp�=q��n><�����
\o�v65�P���3��^��Y������D'?�6������{�&��QF��46'ԭr��㉸�FƳ��*���$���h�"�I�y���J$N��_(tE��}d+��j&������p=�������$kh���*F\�U��-H��L}`7{�2i����b�i�.	E��:�����g�`_�Qq$6{�E��aٛ�ڌ��c�?��U��}�\B:t=��y��
���&��2k>MW��u��b�,�e��
�q�bNJ�?ڊ��0�m��f�B&��orEt��V����z�ФE �軿��cf܃���vZ\Bu�ś L��{�P=w-+��u�/{�'�5�D l��Ԏ�'i*��_�e4��Q�|�)w���0G�/�?f��t���6�t���(�S���ݖ��10�����̾qMგ�$'�l=��A���E�N��� �(�����-����d����;u������������d���"�4��MB�u�(r�k�L������/�4+�v4���%C��[��]�����%�։'�F/�|��YK�\W���(q-�G@��	%�?���W�l��l�����j�k�E���P�ׇt�������q&'ިQ��<$�utO�S���N����R�hZ��"�)�� ���g)���9�m#��{
9=���ǎ��;��X5vu덋0Gg�S�D<c	�OA��FcӓN�@��t�n�LN'�*
k����&�T��!�̾��*���E�����t5�.�d�~��M�XF�FS��>���Z
��
^R�?���ϵt�c�C�z�e�Tٌ��`_	�+W �l�.v`�ح$���)�y�l/7��0��QN&��PX�!��p4�Fj6	� ba>�V��(B6��G5�P��a[{n�{7e����H��`%҂����;�W�uA�t�Ed-���J�"���f��(lvI�2�I�	���ޤ�Ϫd��l���
�{��(�d�����H9bÕ�PHօ������B"n�!*�$M(���ŏƨ�$e�&g�<�1b��rk^"�:�Bׯ�25漣]LC��,�c~
��kW��0�LG$�XP�����|/�^"8�X�x'���XA������
��w�JI[���5x5�)nL�I[#����o�w�;^L	@z@���oF_��>9z�q��U�2���o��q&&�޽�]�c�6aII�����8O����v;J&"�'��̰�ug����M�Hl�F̃�`���h�-ꮗ �K�,�~Y�p���X�C�!0�m��M$K��XI�o�x�g<�(�\pY�䌯&�G{`���6Zg��@��~��m��ֶ۲�$�Oډ	%妖+S2�DًOG�P~G��K8���*���7�o�߿S�$w._ӗje��zX�� �����<4�M�hj;���[��CYQ4{����[�~8�#�Q�>+2�w��m�Jr��^C�N�9���dA���kT8�z�w��@�k�	�?A�
bin��	�V)5+#�ӭ��,{�%�8}�c�S.bXtM^�֋7g�r�?V���~%�.Y�� �E�>�`V��.���U>��(������$� ��є����3��_;�$��7�oAZ�m����(p���.1�%�TR��B�\]cZ�Ө�������ci��'��H��*�q�bu��?<2�Y{Պ�(�����lB�X��CG`^�_��h�h-$�/ũ_3��5\UM�0����1�}��7Dz����H�=�J�Ī��F����R&A����|ŝ�8��!�h����O�����	#N1�OKp�:^cQ'��K�[t�@I�3l��A�#����C��خ��~�����.#R�٪��ͦ��^���T�EG�[��d�7��I��!�$Gg��.�{� &���\4����O%�5L����d��O��Z��O�W���*�J M��W��o1OFKܗ�v��S��7J��UH���W�ެ{}D_�z��SlW�K��rCmP��m%H�m���0�֖�4~�Ǩ<���
���8T�SUӹ��n��[
Y�9���h�]kյ�얍:y�\T�s�Z�)�C�Ȧ�`��������� M�Iw�֓�%`�!�o�H*�G$����5�Ȗ��w�!�����)3fw��۫�����@K�2j���}��d�1\���U�I�I +|G�')�O����̤s,o��TN!�:[|E��_�`B�� B ��r&w_��#�>T�I�F;+,!U!k�X�Xc@��H�5��K���͔3'~DU�|���-�bȬOY�wakk���0/}zů.�R�@��煨�j�ZtS|�d�\I8R4|�L�=4m����H�J)�9�6�d_j��f��A�e��ZA1�2�ױ�� P��,�rkt�C j6�5?��N����g��U�BĢϏ�f���Rq'�����L��b�@����rOw��I��:�$��bFV�_�8��c�lO�@��_���	;����d��R��O�rs�0�g�W܋��X�B�.�H`G$O<�,�����m�S��'N��Y�A�J�;�F��\�{I���c���SV��t^���1��R��h��Q�r��T�k9��Qd��49'o�jK�������ɕ>��t�b�N.��Yys���4Jf+'8��\u�]���
;Q5��w��I�,wo��L@֫!��v�"����}�dlaS"0z��\��Q�5$�GQ����	3���4�B،<�;(6v>�B<w��F�!0�L��iӐ����~��-�M��d��cf�`�3:�R�ߡ��u_�t<�`�%C�2�(E~���A!�j*ւb�0���|����V��%��q�F�=��+Q�pj�Gd��Ɲ�\F�����g^sx��Ns��������D��S�|qKZ��BQ���d�����n���Я��U���ve�{8
�=Qg�naĀ�n�֯�a���f#��l%#z��{������%���#���}6)+�[�&:q��))�6��Eu�n���NL�τ����CQ���$����~�h1oZJ�d��R,1����6����et\�G�A�'��N��G��Ҿq���K����c|g���j���=#� à�a %t��l��'��Jer�eu� '$`�N
���ː(c�6�U)�����6�IC�[D��2-��μ�9&ʱו)*�Z2�))�9�ϙ�.�~���c������.l$�i/����A��I�J ewP��;����C��k:cq�]4�᭶����Y(��h��W�%J�@�ip����[SQ��Ņʴ"P�R:+6�����E�/k��R�i��v� U�;���0#�3,��������ݭ���S�N(�DR�ڐRcXaG�a(P!3"sw;v��+Q�T��Sṭ�x�Q��C�SS�����ˁ�n�]R8.1c�����bt�R��&_�d4/q�=~��m썅���n��{��5@\g)]��A�
��x��ywU&=��z2ؤqv`	9F}���	ל1�-��Ԑ渾�ǖ�(���8�ۭ`/�OC��8R��e�r_��(�m����͡��o$�!���H\*?�i0L,j�w�� 2;r�Ե��r7ȋ\#�v��h��%�U�W��U�w�g���r�o�$.�1�ņ��&=��)a�M�0����gC�Tw��p�3t����͉�p�eG���K���*}�Z%�����ZD���*Ȫ��H�Ew5�

�-�)A���/ėX���(:��w TLu���=��NgS��oě����U�כu$�� rZ���1��ҋPv��%��"���b|8oUƄ�y�o�j�_e����_�6VE���U,GV�_��!��h�����K�w�xD6�p~������I ��3�u��<ԪZE�?ۅ"OS�~�B��a^���'��R!�sQ"*�<|������γ]>Yj��������H���o
Sd���8�\)�X4n�2�s�憫�k^"���I� �\�)��PK�X��	|r�a�ZC�8D��b���>Gq��6����(�/�A.��;b�m��|�K�<l*Ľ۟_z[Z��U�L,��ٺ�f���m�6��DgQ;LIp`r�אV���KƟgs�PM�/Z��B��IGOēEn�#��ޯ��?��e�5Qb����֥� ���� �#�7� h�n?���QC�D�9����S�*���;�q����t+�]
a}ۯ6�E��C�vqn�����8��U���co�P'^��9o�������=��Ļ!9��`�	sy.5��u�f��d�����)e��y�N�f��)~{f���n������֫ D�-1J3e)w/;�(��U�N��;�R�|k�c����BV��o�����e*����,l��s�Q9�,�s��jA%�k��
�9CG�2�i~�6�'fO��k�ԙV7W¼��_�?�\LrG����ɐLH!Z�>�*����ҍ�n�Qf|7P�*��b�ͿnJ�#�G��#A�����o8C�ɨ��RX
)M��ucb8�S����kƬɧ��B��RHz犬�W\����^Ԛ�f�Y]\4���Ұ������Du�MUd���*ֿ����dOM"��S�7&�rő�� ��I>6����$в��0	+.�����l5@�p:>�G�����T��\`_�2��oB֔x� 7�,ݏ$,lg�w���V�[�*��K��fk����*2��B� �;�����L��iS�(�!y�(<Tિ�d>pK,Hi�A�Gu�yEv�L�����4i���S5�(�D���!�������+R��,$,_(>�&2ꉨ�\�.�`�2^����Um�:�[w��U�Ti���
hoJwe��[g��1�Bs	c5��FuLk�cH��m�(�{�r�3i̓�3/�V'�.��<P�ښ�.�=X/2M����/�.b��x�L�����Kf%"�oZ��Ss~�R�C]<<m�hrhy�C�I��#{�)f�Ͷ�l��A�;�P8�`.��S]�G��-�r����e��g��� 37Or�ES�M�L�PQ<�;Z�EÕ.�6�?۝,y���|k�T"Q,d"f�A6c�mW(�U�Ca��Pdw��)�\�+u��5�.���^��w-'W���*(�~sƋ�y�zqL,/�|%����vk3F�e��� �T(	~a��j(�;��8��:����x�dT}°7���{��H���FMu�kK��fc���Ioa<�v��M/�Ç�R:SSZ�����.2&Xѐ�Q��C��;����Q��z�^اp=:��]9�l���������F�?��wnmS{�rԇ4(p���!�;�-�eɾH�->��;NNL�cÈ4s��]ީ�t���ۜ�B3O_߀���Y��p�E4=c�׫�	\Ӕ��A=�}� "�T���هe�8'U���ϢX�[6^/2����'��j�8!| �Yg+c�K��X�oB��)k^��*0��7�:�\z+�Tۗ\���|}E�/}��zìbw���&�q?��AȀ�*3}����'���j���7�F���������vW�mi�4��'���Տe1N�z���e[m���H���9+�(���8B6O���x�P�M7Hn8�5�p����h6l��ŀ�½��L�T����~�G(�D� |<	����8���TF�xA1h����\[�Z�5J��s�R��Mx#�
�����0v�#V�;2��0U(�kə~ѓ"�fOc�<������K%n*_x�B�1�(��ύZf�`^P�24c�H5<��	���oyx��t ��|�жf�#�\zOZ쟄��z<����
�;����݄�{A���>sv\��翇����y��gf�Z[$�R�#��I��� LB� ��+�����B܊ԻE+]���Sa��O���>\��l��J����hp����j^/�����eOOL��%&ֹ�*@��rᚦ�my^q@~�n��a�����0 s��&B^.�hj~�y۾	h�^Z!a�}������}��|��*� ��X�=H*���(g��	q��i˯�i���M����;����X%�7'��\��w�!�¡9�t���1���=`T��9���ΥD��La�i�[��%�~6��I�������3sc6,w�W�����m��v/2$;[�'���J������X$�(_)IiqR�ת�ǧ0��9@v��M5zRZ�� ����ʖ��T��ҰԵ:(�� ���(kj��2U�m�L���`����t�\)ub{��i�3����4�@'���H4:���IQ��A�'����аu��1�|$Fh��ZX,d�������iޘ���V���A'�q�.��xh��ث�[�M{za��	��W�q"�D����[��d2OC��*� ���S�
a</�P�J(�; }!=�hR���*�Z���Uԅ��
�!��1��,�g�4��9�v�)�sL�zU��R�н��r���Ze(����E��Xc'_?X�O��u>��}�Z^t�u�O[0z���#��\05Dy�"�
C5<�EK�ҡL0�M.~�ʾ90�ָ��T~
-g5ȮcC���[t�J(��SI��0�j������!Y9�P)�A�	I���Og=�ly���u9��$�(�x��F&�����n��xx���cm��X2��]�`�~�hv�\��WS�ϲ�M}��:���	�G�[�jeE7O/4:T��A�&z{Z��|@��y�Y8�Ѡ��2����(ª^7����Km��/����Rr��d%�:�?�'�:��xL�����sy*8����0��7�+!f>��ѽF�ٳ��Erʥ��;�)�n���;2#MHAD�B���>Jcf�X�f?�. ��^��."1A�ǯ��}^���V�]����J�x �T�
��CVd��a�L��E�IZǓ|���� *q��"�����Tb�	S)�5�\^T����!]��5�9s�mb�c��,�<Sx��V�T��:CP���}ԈOC �S�=�?S�݁N�8ɫ4�����Uy��.���՗{��9٬�s�j��\��x���6z3;��و�,�P�0�%�)��m��dX�oZ�#��o!B�y���=�^��-��d~��?�Gٵ�?*V�IZ�2�э��z�i!�(A�s�������L�\����kJy��11�� �iN��~��`�ߑ��3���u�"���CD��T�S��fY1�z���F�E[_{}�ݹ���[� X�+R��Vբ*}.Dla���3��@~��L�k]/�;qS:��kte�)Q),��BI�Y��}��3�]�=m�Ö�����si�0�?��i*xq�QQ���Ϭ^d�B��4u�ݤ&��S�y�4����҅��@y���X��5s��\Ƶ�T]S�x�΄�kc��)���\Y�:�#&\�. W��K� S��=�)�>�Q�L��у�P��i��8rp�;���:GnJ�N�AF�J����]�LaP���M�,܆�E]���T	����m�r�|-z�E�)�.Tu�/Z�e�R��o�����N�emG!ƶTW��i�)����׳��z��N[8[G
�GoW���*:G##����olA&hsj��+���:SV!\��اe�#4�������X���������rG�ᔉ"G��B�L7O����18	`�N��%O�ӏ�;��([�(�:Q�� e���
�]ֿe�58d�a���9���;N!�<�#h�S���Hy���j�v|����(p��{��BW̞�=��R��&�T#��ǼCw�b��:����7���N,iF�7�`^��H���K���e�&xII%��]���������7�g �I��P��7��˾�:��зv�x4�A�l�w��h��ޜ(��@�����h�f���)
M�s%��9�ᅪ��qM)�ĢZzE�א��9�&`�� � X4U��\�F�5� ������i`Gh�C��˝S�,[���cv�]}�W_��k���E��w�_��d��#��[y��J�]��Z���7����11#`�՞:/ue�������3c`����$�6N�#y���(*\�s���{�}1-�U.5�1Jš�F���U�5q�� �{$�%�4�aA�-NւH;Xg^�y�8GY95^��A��'�D�1]��ݱK������������#(;,�7�}0sp�R�h4*�tw-[e���Y��m���4��,�q�cCP����'�6��|��09O_y�at1�ׯZ�Fȏ�@�}U��C`�����%�!ۓ�yƖ���C��Y��l߭�V���_�o_�`��VȐ������5ş^,7v����<#�����P�d��\S��\�Zg�BW����e���Q�d߆�[���\K
�O��0Պ}nB����S��8D��M�G��� �<�� ��\�<󗘖�U��C�z_��l�m��}u�t@��c��w�49�\��W�9�((!>��0ף�s�,Եqـ�6��8�O%��Gi���q6�y���'l��[�I3�v?�z��Tz��b�60�U���Lb�ǵ�/&
V	��Z��j���n��X-3�\�<A�G��?���r"�M��g	�)pW�1�&��%#
��Ty�f��tf4�ߠa�@�҃o���cRE���iIf�1�x�6@ �#^�[3<�̪�!��Q�<�׉�"���=M����T��ȖآKx��o13�l���# B��N�c���|Whj�掭��<r׵T�G�f~����_��I��~Fi.X��88����@��?��h���ٴ\&�:w��#/V�ŋ�x{�3���9?[q@�Q9-��C
G>E�U)=z��(ژ�����JP�uf���q���Ob
%���W���v�l$����)���L�J5mű��s�>c��M-^����z�MB�'����������˭�]@[^"ԭ�Zm!N��H�Iܗ�0�<���t�^(���5S���F)��Q�F���/bˍm�`C��>$e!�$(Ϳ�Kv�>�k�!�d�V��j���&�"Ҥ o#���{�.��O�f�(P*��v�ݨM��H����>��c��X�Ƌ敻�Ge����g�ؿy�Gk�����Ұg�z���i_��Všnu7�%��z�x�q��z�bjK�+G�����^�㓍���xO�H-�y���s��a����V^�≏2��]�|r��.�lދ[��.��źY<���y�l�q[����>�M��' 2'���������ܜ`�QWAN=�/���Ǚ7��GC�F��i?7sZ���]9/�0����)�G���진A��Sh߭㋌�!y3����Bq�fEHj����w:T����
bo��c�q�+R��-;o��T��Ot�\���[���<U������D5�_-��9�E���੾,�=4����H�ʖ���-�}VI`H����,�䯾X�kP�l�x�!�j��o�h�V�xW����Ӑ����D�ǩHz��!��ʽ�\vF���6��Tg��M�����N��N;+�C�慑�2�[k���Xo��)=1a<���Sh;����A ��ǚ��䚠�Ew��φKI=���y��u��h X�(��
�k�{�3�:�?�r�ְ=�Ų��Xt��
�&�/UD#�R�S�����K����y�Dx�y{fd/MT�R�����4X掷�^�<A'(�K�Js�{��"[�C-�2��O���AR��ַ�]�YMBdƠ�~����ό�	t��u:c�j��i�.qe��B�r����H��-�nV��Q�M��E��j�EN��8tڻO^��������Fr=��z�*��ѧ�6�����=5�<�D��_�>�*z��~^�7?����U�!�t,C���~�;E��@p�A���oN��IC[����Χ��o�f��F�Ê�uߐ0��4��{o6�����|�`�v�i��j8�\����G��QY`Z�)�٢"�C�lv��}ׁ[�C��s(Pi&�H@�,���:�fU&a��p��Sb�
a�x�<�R��ͯ��t�������{�ao�U����#�����?�"��щ��!���E&��:�7]m��L	��Pb�P�
oB��4'��dֹZ����o��"���̎�%�k'Q���hݙ�6�pQ�fRh�~��+M�p��oQ��8��&RO�y�Q|+( i�x���m{ʝ��醷�?}
�ś��.gR��g�V��M���"�t7'"n���+�Dp������h2�����5j3�X��#�`�r/}��D 2x2X�Mg&-ջ�~�e������6=%��NKE�e�#�F��~�Rv��\т�SVN�#�10�x�ֹB�E#���5Pu5�KW��w�kO�*�i'87	Y��?W��Q�}x:2�1G�p�����S��8��M��Y�k"�J)͵$q�[<Gn�c�i����M')j3��I�J�����W\�K(�L�+O�ǃ�0�Y�����\KpH%a�\�q�8t��&���X�˖E5�]t;qՐNf�@#�Q�tA�Qe�H�R�d�� �X��K���#�[�-��M�+�=�ջ��%�P��2������*P��aU�k��X����w��ɓ)�3*�2a���p�X� [�y����4;J��؝����/�|Y�0��S�2p=���G�c�L?x�_���\=?#{-5F�(IQis��Sh��B�L�R��=����2^N)<$dK���:�:�������Cjޫ� V?ݚVն\��-�B}n!l��c�2��|��@0y%Ւ�p�y�һ`�U�$��� �Nf㇗��۹�μ��EO���p�ͪ��U����Z�����'m���P]��iu��Ȏ��A�i/��(�(A]Yy#:�F}q�/�;�g��Ծ���b�7�����]���MGcNh���A��1��*����,�׵#	E�(++�9�>���	�ykx�u�D�w�-�N����a�s
9Eǁ\F��`vj���
Z ,F�n���GƪQmJM�棽N��0s:
x�N2���ޅ���q:bA����)�
]�B�һڎT�v�LD>@!� ��o�4N^���zLb-�ҟ��:��a��,D�.�$�Z���63u�"�@�HZ\�q���T0s|0R�^>�k�&��1wq(�I���3^�����q��՗�}j]?(Q�Av\Y�Z�0���?o"� ���⟦[�zٍ���OK���w^�Z,��%s4�� =��DM�O~�\��C3���\8wx�?
�m�!JP{"�g���]`[m7����K���zњ{����F�of��~�Gv�K�!۾. �{�����/+�sS�c�D��5@��B	���\G0���o��`1��i%q)�TrHY����4/Ωj�q�{~Ų�\��00����>k�������ԣp����p�Ӌ8:�t��)��]�@�C=�Ե0^lz,���Z0�HS�#���9ĝX�K�6����mT��0��:[����cӘ}�m���P��ؽ��@ɽ�ƪ<��3p��:�L0�.�R��z�k,�S�pw�����{�Jܹ�s�_ɵr�U�rWSc�M9���d2c��T��4*+���Õ�3N� ��*��Ηg1����y��L[@Q��(�fj;�Ni�ʈ5�&�5�dJ'��g<��vj�&��V}Aa�p���V��~��'�&dUj�"3��� �kW�oil���-s
,PM��Y��#��REGII�.�8�ҋ���*<���6g�T����#_�sea퉘Q�k2jCO ,��ע�3m��l*غ��q��/eO���Ky��Oj냇�2�^����W�;��q��M�l`5��ղl�s�1d��o�dàͨJsكz{7��n��[�jQ�ڭ-��n�(����K�\�le��drU%�cѭ�yNd��+_ǚn��6��P&�c�N��;��8��0��'!k��Qc��gW9C|���;��a��70��dς��>���@x�xؠy�K��YuE�A�@ ��i�s�E,m���_t����,�1�t|�0l��Mtp�On5�|G"�s���h�C b'=�,��-�m�.�-U�7�2�9o�(�^ s�G����i�=<�M���w�Q�g;����U��
�YG�k�z4:P�U<�yW�n�~��Ǩ >Av �?�rmռ�)M.J,����9u�I���O���YpN�	/�&<N��Bl(r(Ӎ%��%�vؕ��(�{m�h����^�n�Z�c�"]�zp)5�4^����G2l&�EgM�!���t8�o��òj�����b�"�O�P���a����d��3���'@>����{"g�jH�d��<�)�Yh-Nlwˢ`��Ga\���A�����<�N�4��Q�"dI�E��ȢN.*i�w�r?}I��?��.�(L��v�K���mk����d+�gȳ��AE�0zkF��!~�H�s�C�I1���$��<%H�{��G+'��J�����������Y��`Qת���p�`��̸�Om�U��ܗ�򻙚��j?�B�1����i/��aڥB$OF�Q�m�cωi u�s�4���f�iv��� Vn<��ϸ�侰��S탡U�j�v�}Ɯa���v\H�&��:������s�1�7�m5DCk�'��p���.��#����^�ݧk�Lg`�x�Ǳ����@m�E��%����ҫ��U.t��N����1o���x)�[2���cg@]h�ݨ����'򆦆c-�i7�O[�w6�I���<����F��0w�V2o��~R,D-��ۈז�ZwZ�Ɲ�����C�ԤJ��u�^b��y��������mXS(E����_����b�w��R9õ�;���JzٝGotl�#���X��e4����E���w�v?�w��M
�ڝ)A�*��l�{��)�����ą<cX��)ny����W���.�gv��1ȕ�h`��_/p�^Rݾ�AdlJ%�q�=�w@���yz�I�Pq���?�7� f8&6v
�o�Cņ����y��5/��Z����>��c�\z�[1ԣ�r���7�4�ň
��VS;�1��6QS2�6E���@Ohω���=����{L7���,FmH �F��t=���x��AF���e�
��#ĳ&x�}�	s��ИMi6���Xh=.��	Ix�ڱ�-�E�+�a���]œ���g(��O�ӗ0����%p��
n��7 �gՀ�#��Elh��"����Un=�
,𢑎���x�m���i��B}o	������V
b�J�߿^��c�SAj�E0��x�����FK�t�C�5Y��Z�粭�BPx@i���6�@��J�yr<P���S���G�Xo::kjx�:fGE/���������*f���$I��z>��GR:'*_7�?64�snb��p$�Ѧ����ܰ��Q�c�i��!A�F��l��iEۀ�҅��ל�h�z
�We�r7�V�d����Q���lm� �x�I�l*g���b�_����0�
^d�����*����D�b����zH��U�:�c�����7=S}&t�0��Fb��\�]Co�U��S�r�	w�� � Z�ގyd@tj�<�Hgxu�2r�,r�6�-TaH��F�����U�o���Ӟ:-J��$��?���(�UԌ�s&�?�ܧ+{~��`�y�j /��~u	�����W�ZQ��7�h h�/@A9\�@m�� ����Jf�E ����<�l��f�{?�T��&�%>�����jk��K�#��Ҋ�ن)��>��Rn 	����(�\��h"*�ڽ�'M=�U�^@˭K
��y��O�n��)6]g�}�j�؉U��r��wbjZ�w���U��?(���wJ ,;K�r��q�hs\=�Dϟ��G�ЊTV@H[��{[��`�˫Lh�:y��o�T%��Y*�GI��J�d�������<y��ҩ��!�%��>϶����x��2� O�O1��Do�3_���u��������R�3��0�̌c�Բ�4D��1��J���r����$�K>y(4�Dm:� ��:������G�zNK�,� o/'$G��������ޗԋ���D:�B��c�wi�(��M�;c0�!��E��n9�{!#_|8�q��\̑4l�<�<��I�U�A�k��g{RA��<�'a�*�d͗M�C�p[.�мw��)�S��
ǯ-BJD-4.3�A+cL$��S�XE��D��]��C-&��F��-�Hܛ[ы�ap�ZF�����zmSuＷ՜F}����Du��q�&��M��Ѯ��vwX�㨰K�Q/���hZJW&%�d|̤Y�מ�ܦ���Ya���'lq)r"�k�
�Np䒓�S�HK�"�����61��]L�/t���YE^Y���ş��뫑0*��l�+jl��q�� ����^�/���8���'������M���i���8�x=�ĒC�C��}�p��硠s�Z<�~����;��>S�7�
X��Q��rXpGo��`>�ŀ�N���I�m7�Z�?��~�"�l���^ų���4
��E,�����I�����汄�5I��E77�x��&��<W�c�uӆ���|�E�|���O#��}�e��PG�߂�y�I ��J���ʒ�(����z����Cy` �(�)��lq' ^�U�V�P�Zi����)�~e��ƌ֍_��з?jQ�A�# �����&����z�ž/�u}[��Y��̆�DIz?����B3��I��Zx����ӨON|��Į����m���)r���a�ſ
�6��F����������?��0�('	*֒ņi�J1�@��){�,&߾j�	���a�!.,��|�]���(e>Eվm*�l<V|�XV�
�tvo�[y
w���i�究�������Q�B�&���u���i{b0����� �㊘�����Li��m�W6Vt�����-b�Q�3c����u?��B�%l�OG�}�l�w7���c��|-�+��:���e4����m�E`�]I�qa�df7�$��K{�[�:_�SC1xa�����g�[�������(f}3��mK��3���-L ��C��ji1%'p�:L�8[� +�g�>��T�s�0����)
�/2@x���[��y�_�� X�����Q�#ֈ�, �'���A㫽|���#�@/�]�B`��v�rC	jW��:RyO���=/�tb��,l�-��� �mW}ȩ�(f!P���Zq`���u%�m�����-�Ŀc��u��:(�cw\��ah��F�q��83kL e����I��|��������>���}$���t$�.��܅P��4�0�,���]*�ܘ�����V�+VU3�Mů{䎋�����A��![3kNQiy�QdhK�wO/xƐk]ۇ�'�����2�Li�"7����+��+�d�����D|��Pn�mv6t�19)�˳���h�T1!,�Շ:. ��h>ح�b/t�y����:��g9�t�Z͹g
}�Zm��4� �}[��F���ٻ��C9�2�a�l��ʴZ��R(�5�h�F�	R�I���y˜өf'���5 ӽll(�nk�z��zQ�bl1T��|��6C�)X�b���жN��/[��FZ
��q�F�~+`1{U�HA��_���Z���jͳ��O�t�,���*�����v�4i-��fj�z�D�:��h%�f�<;Rނ,�2̱W}�6�.�o��H�������g�0>��얇j��=����-��7N�4�3-�l��E� !���ֆ�߸	����(N�j��N$^�T�sf�R1k�TQe䳊zE��m��B]{�k`����z�9+�*���j�P٦�n�ż�J~�2`.���w��#�%ְ��rYW�ӣ��:���A&�f�
¼�&�B����)���w`VV�`WP��40IW�����+H��áp��S�:&�4��xߦ%u����8x(���C^��CɷӬ�]���a&*(ؖ��b9�X��=�/aթ�e�|m�ЮI� (sB��KjR�� ��2�o�Ʊ�q�@��2I�i}ji9�oT�(܁w;]Y��9���ZEK<����a>��ݨ�h��[os�V�~�Ȧ��r����^h"����_Q �A;�b�b�& �w|@�]~"���x"�(�oΝ���=��F��G��{![A�X��@�0D�X��2G9�m���ܶ��J�W���.`�~Oa� i��?!*�%;��bz�/!���+��\ L9���A֖W�b�"��Q��x�6�/��v�m��@��Z	�j�R�{�W�'k-xl��mUGD��y�������#�]�:Z��B�P�C�	؆ ��k�z��:[,�418~ϛ߸���j�g�l��UG���%$)<�|@k}�޶�<�p �&�\��4��7ë�k���ޛ(��4�]jbp}Pf�E�B�h���d��
��f���p�&(��t�K�@_���6
����NJ���w��o5���>#���椱|�p3H�W.�z�7�n8�M��\��-ZT �^~��Cm՘�y���C����,�6��p�5��|<������� F����N�V+�C�l}���e�4%_ N���7�l�:��??5�VT��ƒ�T%�lo�!�z����3	:=��n�q�mT�N����y��42H�$^-p��PzϮW;��⼒�qiޱ����14I'������������	p�w�K��Ex���B��`cU�֛���q�pwL�f�t���,-/�ɛ���F�u�(ؐM���="�ؾ�hYt�Y^sHM[:��XU�q
�<	������ݾ�����	�n����s�(Ԝ�\K��M6o> ���כt��n��<�v��o�6<uw?^`=iM�Ӽ<OcW�}i�ү�1n\�k��-z���7�0��T��]��V�8��E�����>X�����JW�7bF3����]��H��>�m`m;r�1�Ж']S#��\�f�.��{�D�:�X��,���ӌ�!%vQ/����.S�&&�5�����1K$���:��=
lU���.i؊�I��g��1�����!����PU���0������}	c{ڊ� ;=�L�%ύљz)\�u�r�n �����f�w�e��K�7��o�_�Z/�Ψ�)N�Z� D�P����=�/{������>���Z�4_�W(�xX9�� ��8��U	#�۶��@[b��,�G���D���(�4�bT~��(¬���I�̗=G���J�/�� �x�i�����}z�#�E��
��ʮ�P.�1[�8U�O��w�D�2J�,[P\�k|���O�Qu����J�T��ⳗ��ES&�Q����T��EW*t$ c{�F�	��,*��wV�vW��KHDA慽�.~�%)�����0$#_)�f7��iM�����ӛ-�ә@��"MِLc{�߆�]���_4Iv�D�/��﫱	�TZ�!u�����5�#]��"��'�=�M"7_[R$1oE!ͷ34�p���琄��i.���oj�����X�M{Ps�%v��$��M��y! ����h��!_odnI�v��Y�+�>ov�MǤ��.
Z���ۄ5���~��It�j�]1��SDف�^�N�4��ͨX�G�I�S�gk��ܤ�K�	5Lx�ޙ��ގzUp5��,�e/�3`���WAr�������<c+tΤ���9�?!Pv�� �v�(xa_s�6� h ^��>C��!IC$��C]8���6"+��-_��/Wi�� ���)�m�ap�������y�I޲�ݭv�F�Ƒ;1��h�!ވѹ'����+Q�G1�R�;�iմZ=�c,�M��pKdo�<q��?S�>�e��=hQ+kr���Q#p�&f.`5�M���bz=�\��9٨���%�Eh���i|hs�Y�Z�3)g+��̞ !4
�W��O�:J6�2;�����͞:���XE�A6��A��F�^���Z�һF�����Ui�Mq�^��x�'��~8;oC�^ħ��9��z1�m9�@_3�ҩ^��ġ�_�5D�*�fN�r#e�M�g���G�z7qdO�qM�y�T���lէ�'������f��V�I<C
��Z":ᇋf"�t�L�����"��AfZ��Z����۝q��ė:���-��������H���A�Յ�����L�i��ݶʇ���/z�^��Vp��O�&��9��X�����JAF.�7i��7�|�����#�7�ɾ�������vU2�+P+AC�o�A|�1n,t5{�t����u�d����O���sɬ\*DM͎�{�o��s.4� ���c� O�m��$�����{�bN#a��Fك�?^ �Sb�z�`�tx�N�N|Y����i3�����#��T��c��4�_�T�� <�%'J/έeb#?E�`x���֌;u-�G�H����>��|��=Q�8A��t�DWe���s�
Nńv���7�r�U�H���+j�������*'�0SByU�-$���LT�~�k�R�e���߭X=et�b�3��1-%ay�?{��5�X��ȁ����v~�'��j5��Z$�B��v�MU&?Y��@��P����I>��]b��}tn.���6T�u��Q+K��Æm`s!� ��턲MQ��,Ix7�հ�1�H2�N/[�A����1��5�!y��z	�>��������my`܋ui�V��oF��E�`ޟ���Ƕ6rڶs��1����ƹ�{� +;Q���3H�1D����X��q�xW��S�?�.�*�+��oJfc�|��t����a�6U$k�ϝ�QxjjUB�#����9i<N�v��M�ЛȀr�i�!	���z.�E����#�pE�������w+B`ң�#��{x%4\�9�a�F_�s��r�\��%z�ݨl�6ڸ4���,ּe�&�4g���!湢x��M�8�?#�a/e�h� k�����K�s�J�h��4�-��.�-Y
�x:d�����f!��*>S������Dr%�#���	�i��[}�P5�Y�-��t�w����R�k�5q�^:�4]�<#��l��z(�-[¨k,Օ5�T�c �&$<�V��eՌe��&eR�k����cK��ձĦ %�Er��]	�5�{(��s���s[�\����c���#�5��,1]o ����nx���qN<&�����Bv;�4K����b:���z����A�٣��!,�?�����;/3ר���z(	Sq��QqR��Ok*��;����9A�e~9˃=_'�� �Ym�E�����h"$�[�~�}q�y5}��|l��a��0D�)縆:�hB�ŝw��Iܡ|Н�9�6_����R�v��1��hҽ�' 𜜡1!���(^@aF֐������v]{��t,��:m�5iIR����}},��C�����81��,������)sĻ%]�3a3*��Ѻ�JnIH�Rh�zs_��n�X@��&^%O�O�ک�Ҧ���Ê��Ǻ7 �(S��_�G�"j:=ي*�2p��4�h-7k�3�����@�d��>i�]i�e�'������QL�7Υ�+e=�.�����nX2��s�������!�V�q/XY
7�. xE.�O��u�0���U�t�R� x����Y�]]�kI�G�p��z"K�;jz�֓����O�S�;m/-*�֑��ܖ>����]�X �r�r�{I+߳f�b��(�-��I����ݹO�Q	���� 6B{%|��  U�s�/p�;|;���th<����+�wU��]���������uC�iF,Yi��_�����&|R��۞g���̊þY~�r��"~*�E�R~���<�6�In�݄�d���?O�}��5M�Y'�X0��1�x�ygl#�+���xa�u�4������^��Jo`^(��쀙"��X8X��s�+�@��g���a;��1J{��L�N�.�1t�K1:4�
�Oj<����n�K���^���1�<�Dr���a(/|���yW'�J�̼�c��E��(�.��X�;�k�S� vu��7�w��VJ��Q���5�G���ޑ�?<�1^ફ��)g���*�D9E���Z�ۛF�0��U>h�뿱�y���L|y�劓n@u�^�3�ƭE�����|Sz�j=#.��qk���ӣ�D�sD�8~�(3�'��+�e�9�ov��k앤<1�}�0�HCg(�[��1���gOB���Ѹ%�f��jpP����T����{��[B��-��U�sb���_�VXE����1��O��Ceg��53�r����RЉg����ƈ5L�6��K�`��<n��P]F=�����y	�}���Gm���x��n�j	�X��DSk0�O3��|v�q�5s�Vm�B���]7�ÿ:q�`��X�q��:���|�[�w�Zn�0�����	���=Y�׋���|w܈Z���q�[����dk�}�vsV�l�M��ux;����W$�{��`��� �W�!\Y3��C�x����r�ΗL���pw.E<��-N���C�а�T�NQ��z딙/�<�O`���Z�BV{�]�N���O�ݽ��F���W;^|�P�2��6�1~	9���Z!�1�M�s�cv��n��Z�.��2P]�n�<�R@�g
2?3����2�|�{h�>
�t� ��꽟dR��Ryf|�DD�l���@.X�T�;W'��P���=�^�/��-�������h��b�+���Q��D���߃���s���RwNm�$���J;�ʳ_�e�:z�aO|���@���1gN�� ��k�t����|d�Z`�q ��
Pݒ�Đ�h�۫!�	���rS�������M��$(��W7�*hF[ґ���"�IM��]�ֈ�Q��=��3S��~z /=��|W 4X�q�%
锔�B��f���oJ�C�SP�|j���}POZ 6֩Me��? t`"�94�,�~�U�Gz�c ��ű#�F���7�����Vܐ��G;�l��ő�T��X��d�3,L��Sau@k��jx37��w��cQP�d֗܆e��)��"	�4U��%��c}�Ʒɬ���M'�Z���j�F`ءB[�@�_[ʮ���D��]k��$�6�\��׺T���q��+��0��=z!X'H>9�_쏤@oɉ�>'��J$�/��-5�_�V͋��Ƒ��W�K+l�����?�.K��ՒHr]�אն�洕Ω�d8�����Ǣ4��K,���@+���k�N��u���C�Ye�e#�q^�ȣ��љ5,Djբ7\x��7jZ�s4ק��]��j�ʹ�1;�F�Z�R	,��S-�4�y���-���0:v���V�_^0�������4g)�Oߊ_ҙSK\IcSw)X}�$�J��>�/at;�KA载�w����K5�/�N�+8P��$w�-H`���$F�]@GqңO�H	bw0��l�XZ�Ő�i/I> b�v�����ĒR�<����8a"��r	�C���<��X���J����94T�?2�M$7�����$D᪇���9����m+����c�ն��>Ct�˚]X��v7i;'p �V�0��P��i/Z!�s�; -�7�(�e6�|.��5�UAy�c	Hc{�"\�,	;��q(Ua5��J��r�<�AĬ�=`�V�����9o��J�	������C
T�Ȭ��.K������p��/kw����M�����m�kkE�{xfd��X���ڦ��)��`bh���6�a�x���'�rP5�D��d�'P����7��<s���ð	�So�C�܌�V]����{Ts��;����#��DQ���n���4�n.�l:?���
�&�`�Q��ذn���#g��t���7ߨK���o��,z��QS���F��@��TKI� zTo�����6S�%��d鞐ZL_���ǫW7n[�[	r��%4��-{�M��-JC�F��lޕ�wK�ι��3�@�x�P�@���Þ ��l�e����ZGt�,��Y����7��!��3��*�����S��Dx��ؘK����I�Fk*�[Y�� `����A,��W��;́�IvDə�A��c�>P�Um�ުoZ�-���l*�X��?{��/�JZ������T��]"�e'f��koO�˝g+k|�A�GV��Gh�\A�(V{�pj|:Ѷ<����1����e8��״���昇�x�J2�5ڔ�RO���5Q�r|:<�t� I4���Tg�[r1�c�:�2�Y�N%3��i,&���"��njR���z&�/ǰ1��̩袃�j�Nq�"�u�T޻�Z����D-/� �ose� ��Ɲ?�^m�9�k	(��GBқ��'4{Cr��񰆎���</9r�p�������u�w0t��\��EP��d�U�2�	��^	�4&�Z��'$�i���]E� [0!2Z0��!L}D�n�Kp�T�Mr���{j�D7L,��|9���觕�=�ajx�7�^���T�
P�LA���#&�;��O�v7ԧ/����|`�5���՚gQR�X�.x��N{#�
���h�c1T�D�A���t�v����� �t�|�Ǽ/.t�5!U0���[vu��]���Y9T}J�ѱT�����>��4���N�E����,�q�����7���<e�Wg�f�c��Ig�~K�Dii��|@C�l��\³t�.;��\7�XP��J1p�ThYǫP�4w%v^�d���N�_�[E�:���:�-|#�+pm�.�x��]���	`�2�*~�`��{N�$g��)�0o��� 5�3��h>L�vi�2��ÊY�N(�Pv_|��,h3e�lb�D�W�&���)���o����1/��L?�����1ힾ�~qe5���XTE�
��: bH�BD��51���fO��N�(���A5�2O����U�VOq�T��^sX���rDu T�!��M�)j��3��7R^�'��$?��:��q�yA�>�K��`�'�еմ�C���m���i�=ElQb��\\SBC�~ZuvX%YJ��T���Zm���:��b����'������9�k���p��xIǷʪ���J�@5��+���%�R�"1vIޞ.EdN��s���t8�����K�;粣iHŘ����D�.l>,)��>�q���$���k+���|2�V6�4y�1��8.��5�uN�yf��0لU��_Rg���f�;�s/�/�?@�f�.9C����G��D�y���,N=�B������G�����p٧�<��ۋ��9lP0M��T:�A�B����8z��¤j�yE�=s�ѤC0`�V�_���s�	����A,5"֖�n;?I��.S�$.T�QdanCi &�j%msFw���F5ѕ��0�#}~a�UHض{N�!/}a���J%&������JW��v�۴�<���\���r{\��y	��d������5�����8B�!�tt�k���n܍w:�;A�09=h��,�������������*��߷L�ƾ��^�ݠwMO}\"��O�ã��tj��I���Н-�*�i��s��'����#�  Ζ31%MpS�e�0�f>l	L1؁r�A��	kEo�����U�����L�u��S7�JDd!*�@�!4���M{�%��z�K����{H�yv2T�����ʐ-�)X���L<���I�p{��}C(���)M�M�1��I�NR[iY� 
`�����^������JD�9Ò�	��ؠ�fXX+iT=&1��fߣ��wZ�a��X�fi��"���=C��+�{Uh�/����MR���(��?l%���C�X#����%~��\�N� ��/5$2�gt3]�Ƿt�=�|Ȳ�L]1y���!����oY�e(�au��od)�v�xw��ަ�T*�x��	`�������gG���D������Ȍ�� l�>�c�L����W*/� :m�Le^C�a����O�s-�j��c�,%�3N���쾛�P�QӨХ�鎭zO6�A�l� ��CX�
�2#1^ 8�n�߽ԙ�0��P�h}Ѕ��[��>$����}��d�hv�-��"�"�m$��|��
3�yn�\`�=Fx��g�˯tF��� ��=�����<9�G׊/&�oj�̫�*�z=�]�{S1��A���`^�&W^i>B�]�.%w	��8�(��QN��h6�г�WL�P��ҽB��>%L�#��!]݈������!Ъ�k����d@�����T]�H�5�������ɜ�rv�+�f�l���cm�<�su�3Ш~��e��=a���S=����u���nLS'Ed���v�QS>��T9�j��	>�4�S�.k8V=����%N�yPcV/YJ=2���ާ賮�H��O�)�����Mw��$�
}q�ݹ�_W*��p���0�@w�Gq�[�b�
��~f�3�&���^qށ]�I��j�Z��y���K�y� }���y�ӂ9G)��Ȼ���jM:�x��8�U��Et��h{�����No�&~�» �P���j��1/�:��Ro�"�v�X�Q5����)��<��p��{�XČ�1m-��U��AP.(w�<��c�d��?0f
����q[�݊q��?��}D%�6�M���b�%̻ƍ�F���yh�vM�R�^���˨6V(�hΉz��sU�Ɨ�3FA+�j$`�V��� x�?#t�4����Ҏ�b�H��� �ڦ�˃}a+�e��Ԛ�q��i�j�k��f�k툽��Ѳ��N5�=m|r���Ǝ�s�A��A��kHM_��������}�8�0���+q��w�O1�·H�k�儷��3	��`F��5
T�5?K:�c�tEC=A$�[q收 �[+
�c|
�f��EB�������w�Zpڍ�f|�>PB�K0��n&_�]W��ĹM�X��5��A�9���J�_U��ȚP����d��~��5�y9���Fb��n��gm:�K�Qߖq��T'��$!T�����0#f@���: ah��@��������/q��ʯ�+����!�EӞ�q/Uo��5z�'ʨ-o�Dk�2�u������tL��^϶�9���^JӚP��#UE�P	�V2?vH��wǧ&Ar(p>�ؙӓo����C�|�M j�$2�͍��z�b��B�>'FN��OZ�g�����-lLDGC9iyѭ��R�	T���ϗ�ZO�&���̬X� �ZY4>!��b&@EYR��"Q��'��?���[�C'J�����ڧ������P���v�Q����ռ>��*�v*�L �7�0g
�4����ߘ���y�U��W�j �9��Im�����!�m�I���#�r��ǅ�,���Y'I��0B�*����fG�5��=��ӟ�a�9�g�#�/�P=��*���Rd�l�#� P�V�t�[̯j�yz~�e>< �;�+@��.8�aM�h����=�N!�����݁���A�L�R�D,�.��U� �ɬ��.=�&�?������l����z�Et�ُ��t�����O����W�W�1|V>�"E�BJ��?sjx��ɔO�ߑ�c�N�9&$cX�<�������ӕ�b���vV ��F�0o�?C]Y/�S�cc{嫓U|�g���Hh�p|�]e��y��}�d��Ϥ4�C���Ń�:��Z�w���䐼�`��Z��C�X���,&�4��^:��Z�}d˕G_���Ke�}��J($�̝�r��)"�ҰF�N,"GP�>j���la,�C�^���I��#����4T�k���?(�C	Fl����l���}^�!rT;eiS�V�Er1��}bٶKdG	�\˧��ms�	M��Is��W܅᭞_14�3�B-9��'��N���k6���NZ�O��l�h���xrӁl�ñx�棉m+ )��6{M���D1�e <G�'��1� F���՗�����4&��'>�����a +nJ�;$.���.���¡A�MuLwG�+��3vb�P,�?���v�5����˃ -�2��L�������%�F���_<B�0ma ��8E�.V/x���0����Wrr������+.uYw�J�R[�&��*����t�ҘDB�c27�X���KY����B�^����ky�}���t�x�w�!����vrJ��Vz��Sx���ظ/�<��0yJ�ܥ�����3� B����9sP�T�%�'�k��"�Y)o �6������ʜCi�Ġ7������_e�U��%4�
f�y��V���s���V�2G(+UB4�
l�=����7h��D#�o�y��9��T]e���҈��LJ��N �_l�,�ί�q���j�����oaa�j�����iv�(���GR�i�y"O���\W�Z)-;�V��9bhkqfA;����r���e;�NW���#���Z>����س"b����ހ�$vq�A���\�re8��_�ǘ��֣��.W�Kh9�[ͦG}VV���t�p�˘gY|�)�t�%F�ɑC!`��Oҕ���0�h���A�6��8�541%'�V(�(pX3���Q���;�`��!�j�����b�N��D{��4���jh��v��b_�SدU�%��9J����t�FB((} \oi 3��������]@�$J�.`?�-�Gr|K��(��J����6<<��8˨�r�t�sND���i��G��0`�X�t�Bz���k C �*-.�R���4����4�jW��UAd���hH܎�%��wܮ��P������ѿol@&��;z��m@ҝ��?��b���:c�=�u��7��6��W�y$�)����a�[;2?A(�<�$7�K��m���yڂ,��x��a�z���k�>[2ڛ�&b��RH&pੑ9Q�R��oo��m0U�T-\�i��o�B�/�{�+�p�_gt���j��ju��USL�I��J�_e�t������ϧ�_b7p�N�4G*�-�2���:l[�_���G$T&ߤ���ڱ[���|	�h`� P ��Jn�Kƻ4��8�0�o6��X�y���z0M�H�#"���>\{L����k�wFE�Ր�M�.9��F�l�wa����汘��:�LN��"v���H�#Z&&`��6� �2�j�Q!i����YW��+��� ��/�*��͜/~��b4ű���~�a�W��c�ˤs�6�����+�ЫYh���K"�_��A{�,��fl)-'a��:�*j0�k��R��o�W�!l�(�� ﺶ�q��տ�ϥ��9O�|=UXu�=m-���SM��8�d�
@��k(*�����Ά��U+�v����])Sش^���Q4�+Ǖ萜��1���ŷ�l�_��j�@Ա22D4�YU���So	���Y�G֘i��������Hp�u3�oA��+ܩ8s���Ά����W� �aWT��3=(�d�90m�]��=��/��hhH�?�5\��r/{���s&�bO����+?���!�:�j[d.j��Ns���.7H���1ΧYr�Y3�ޖ@.z&b(�}Եw��=�\Q( +�s�	H[zJ.���>�����"Z<�kn�J��Fc��i��zڈ����e�+���Ɣ,�/��T���^!�Stg��K.�nR4j�r�ǏT���)�w�lǬ�Q��m����8�^U����ʓo�f��UpCB"�����%�]��oM�߇ f�s��}/��!S5�
��!����o�?:�Ηj(C}m�]ql���|Xp�2��Rd�tEI��|���Avml)��'�.�������<��(?�[{;ݎvX@-�Ǎ�alŶB�����N�}e�?��	I���L�	���rv=�f8�U� �;�]�㳧������`�j��`�SC�'\�7���s���C5�c'�������N�Z(]�{"%���٣)��e��.'��|q�Fz�����3��B<J�#"J_�2�ώ�H}��B�F�i�Z��`Î�'@��,�!�;�'�ot��!Nn;K'��ԛw����r��"�g����
Oi��ƺ�I	��YXW�'!��dN�UI��������������o��+/�Nɢj$�lН��]�H�C���_1�̣��;Kἢ�$�d��1v��0��8x���F#|A��t��f�#,��$hB'��	�k��
3	@��LXWP��Ѿ#�<Tc��W� v�,��!}?23� �t�-�R�rt��X������� ��"� Q�k�����&�9n[��[ɌB��tq�"�g2i����+��fS�o�	�5U���FЯ�^GCbK�s�����.��J,�_l�r.��j�q��.�,�m/s�a����Ѻ�����3k�&�~1� �l "��Vܤ��r�<�����ŋ3���W��ʖ���pgQ	�������M�N�%L�(�cr�^�b`ʠ�OZ�w��B�n���^�X�=����z"�ނʯ&�l�w�xh;�;lQA����E�v��Rj79��§V+�^zj���c:�x��!�7� ���vFi�֘z��W?��ff���^$���al�i',��t2��y����[Pw��N��V	�niT>��A�8O��p����x;z}��V(��e�?C��mS�����>ܣ/c�wU����P�q8�[f9�W�h��MYa�g���N�)`2ooMi��4����8&��cQ�pHQ�/�1��&����8��N6H�V�d?x\�~(H����a����.�b.7b��H�ɀ�v5�j C�� �_��9:����q���A�n%��o��z�H���Ah���Q����M���D����,�aq������Qvũ���+z�p�Ȩ��p��j@�+��V�ޥ������p运|����h�����C4q���ߴ��j
T�*�͝V��4�>��O@���DC�����]#D!_q�����j�]���(Y���x�����v��U���U�V�X��b?����?�ϧtݡ��$�7��iV�Kp9rG��Y��Z{��Z�4�K���0�V(q+��-%G8�(��瘓	���]#	�����r�h��_��'��V7�k��Q�;�N#��%wE�w�9ҏcبT�iѫ������*�0�������6��Hёep����={�@�B,�wp��"�ٵs:k���1�%�!dJ��v��t��HTB.q��ށq6;$PZnӖ�aju�H�@��8gf� �A�������ѹ[����G���dd���]&Tt�R�2p��|��<M�`/a�΢ĆYz�^f�������wR 4�Z����	�{�Z�5[l���LMG{�Kk@��1��F�Y_m|��>�I�0������h������R��`\�?�4�u(�9x������w#!�Ĩ;����?�~M��,j]!���%Y#�f�;'�0.����,G�	z�d����^Ԅ:��2����.�E+(����]c�U	]�������P����D'yu�C:�s'Zaru�b`*�,�$ ����Bm�c��:���ai��E�wY��W�0�w�N2Su~��=ִ%C|�ݚ�v���B;C=#�"A�Uc�,�S����`�k_z±���9wp#~0��w��\�/��@�KW���c!���b�����9�J\�F#\���	�����Ҝ�P~�A��W�C�j�ݘ)2�����w��D�[67ʝ(�8>�)h^ΩeW���Ն��X���|�U:���!��z��V�mM����L����þT�l�')53	w�)S�c�1������:u�!7�cs�A��}���D~�b����4�8%�8x~��B��9������i�S�l��fz5��+xo�!LGa>k��dOץ*,����o"���a1��VV�`���[�Wr��+'�p$������g��	 \��J�v����F�0<o�N�e����4)C��q���[�u ���yK�l��UY����`��;zQ�x.���[uw8M�b���7zI
���m-���T�3�� ':���A&v昑FSr�JE�v�jG�d-,©6�L:�B�m��(Ha��C��P�D��R����_P�ϱ�!:O�|qN,��^��Z"6�Ч�-�z���hKn>���p�_����N�;�e�{~j�hN"73�)f�~�@���n��m��,p{;�Y�����8�rMjAv�D�a�b��Lۀ,B2��]A\��M�#P�vݹ����=�&�3�#X1�|Q�"�s8�,���N\�M�6�:>6�$���H9�Wn\g��Myt3�T���/��4�Y�;������.e1$[�$^P�v���Lj0g�^F�u�o�S�rӾ�����ܯ\.v�=�
�O�zd��>����e?�ֲM�nt,���l%Wn�{���+ϞXoC�m�V�2�5����ܿ�IY�U��|���uLd&��]�lgd�&o_�5�U;A_��W�(]�~��N���xX#V�.���/�Q9��:���S�+��nJ��oBFp��e{b c�� r �5+ʩ�� ��m�Nu��YF��C�.���L��������TB������h���A/H�Tn~M0u@���QCr�>G���X��k��M/����61'�3�i���k3�A����{:�!����oT��yW�Z	a���}C��yp�Fh\z�H�0g�T?Jz�'�s���)2U̅}	U)�����t���} �_pR������ y�m�,z1��M�c�_��w�Ar(��i�~�QcN7�j�t޹a!��g-�1S���V�Gl����T5��[կ�.�i�]��
��5��xm��BB�P��(��ɪ &��Z����@�x�+�`l��6#W�h����'�?f�	T��Ձ8%~����G<���7U��1����^$�S�L!��t�U����!�P��Y�t�d
�0m�����e�(Ν�՘��r�2?�1��q�ۅm��0�����-���\��ј�t:�1���������������@�9���.��7 V6��u�����g)(������}��w>��r�F�uH8IO~Ң��hq�3>�[["�R���zw����� ����_�	Al�R���+�����C���D�gg���Ќ`��`#?(���AxÄ�X��rw��N������̼���}� 5�t�z�2�GM�G}�kB�v�-�_�	�!��vy(��o>�iV�X�2���%�S��κ��,�",AzO*���[H�G�4�>��e�Պn*o�����@��W�k~�lVJ"����J^SY�~�w5�m�MP�޾�O�/ŐQ_�O
8��ҫ �+��Ը��*�A͝�L�np �{DKw��z�g�#��d�ꮽ��)X�nq��Z^B�,Х_0�⑃Խ����l;̏>2� x�e�~��cT{����O ��ɫ~<>hű k[��(o�۲{Ǐ<O��wf���l�N3��A�c�W?� `�T��d����X�;?$*�,�Cr?D�E�(b��\�������,h]Q�����j�S:v�?7q�9K�E�����LN~���>Zc�b��'k �JX��`��V��s(t1�⁝%����o����V���%�*����8�?�Q�.w�:Ͼp�BmG�h]>)3o�ş5P��F6
��.h�b�^�\�ZK�Tc�'�/21s}�
,#�w��S�<�яF��rQ���3Җ���j{
�,O��������V�J@�-
�kw����3(�s�>Y��'��B��k ���m�׶X?��s9�q�]c��5�+�R����B�c&%M1ƒ�?;�!��k@�W�t�n�x�a���8?��M�[�X�_���Ty���p��#w����V�m�_3����������J�A^ᣥ ��O�_�Uh~��S��YvGjV&FQx�5G{�aV�/<�p�������9JZ����`�@��ecTaHn����I��<	�G������Dq�I�����-�E�s����CG6wr0]�����g4jdY}��PU�nƸ��ҟ�qs�!�*G�`9)�~������!j�����z������+Z��FO���Tms���z�΀��),��G�ײ����T&��ᷡ
��GH�p��!��TO�6H����t��%�#ic���;غI=/7�e)S�r��-��v�`B����v���r�ߜ���iA�Ec6~��ożb��a�L����0{z�"��8��^�4�K�P�ʺɌx4��u��罕��a�B_߆8/h��	;M����x٠GM�V�T�m�;�vؖ�m%�H�D:y ��&+��5\�/�f^E��|b=�0���tz�(hy\*#�+��3?
{5�9�y�$����I�.F�'���{n�3�����P]'{,�m���\�������#�C�[�܎����������F�����D�:<8T��ŃJOx�oG8�W:{y�;��2�_XL�N�t��#ݱ7(��x^P�����k:�Z��p��;yYR�m�{0��%$�76o�����͵i�2�ݩ���|�6V�|E	�a;�Hͧ�#�fIB�6��V否��|V�`2u�����1H��р�q@[�u�y2�d����I­����&zk����y����iq�Z��?��Xn�|�y�5���G�+d��WO�:��(�m�����9�yU�1�eg��J�%;@'�`�L�Y������+�>��:#F�Gx�3�,|¸��_��-ە?ϵ�l5L�5Y�d���ߞ�؍��C&x	/pע�$ � ��f��z+�m�Sf���;E��s������xs�4<+
�\C��W�����9�ZJѭI�_g��ƨ�b9����g_ջ�O��ՙ>��p�v�������n�`�E�j_�+�Xj�#���悰�7���1�tP�#tEEo�?�:��v)�׼i�իf�+_)�o��nߪt-��,�A��kʑ��Sh��s�'�Xt�]<K���Q,Y;Z����郮��+�+�h�3�9�T�xM,]ؙ�����:���>ǋ_ �t�vv�Lk"p�jM��H���.�b�p\diivl0aOK�j�T'/�y�*���9�;|XH!����w��B8���Hހ|��j����v��j�6��>��x�lP����LXH`@��������-֥��r2���?�D���K���̋U��|�L����6�j�������֏~�~��ݒm"�w��lu:��AEd����o�I�J�5c�d��*�&�(��D�has����ܨ_ʍ�v�c�cd��P�{_�GCt5\PU�ONDS��jNm4��cZ�#{�������I�(�bO����'�;��y���b_~��v/FW|��j��4O���=�jC�L/��v�9�b��gQ7&u�C�7T�������5�7Df/Y�f�Ϛ��1�)��#q��׳y���IZ�Y�GV�}������5�o(�<����Q��B���P4���P�V���@	$������}���K��@�]�C��bЂ^茜}=�.�bVQ��Mn�w&Z�h0
P6��N�7؄k�`��Q�!)�l4⣅̳�K��iWZļ��g;j�FtZ�N&UScw��<�i^;I���x��i�!jO���Gxt��?odcD3�8���r��-nL�:j��يe�*(��~S�߅�W���!��S�"io�"ƑאD_z9*c��@=�_�Ե�|�9!��������U�@�Z)C�}�m�B��% /����r�+��X�T���!�bd�m���e���ȕAJ|�!ߗ���!��l����|�r��"0J|�1{��9wv	|�l�\��V�� ���jЩ�|ӖX��[�H�����Sh��zFz�"�e^Lk���0�v%����*��=vs���y�㵊���1�$CZ�>����e7ˎU)/�'Ew�"#��](����I�/H[�~��>87���MP��v�bogϟx4|a��>��V����ǚȭ�6�'�M���Jn�w�٤�ކ�|���t�|��!���������A�fm�����(��a��v�]��jŪ���)y�����#�|揟�z&$U���Ѐ�}�E~G�Qg����A8��>�O��hY��QY+��,�&~>6���7Kv��I*�6AU�g�YuW��(��}�;Gmn���N/|x�=5��[%":Q��A��M�+��^	ZL.���L
d/�Z���ȅ��P��i���v<��,�R8�z ��qb�,A���1a�z���T\Wpϴ���r�z�N�]��g�ʜ����^qV`iK�wJ�h����q��_��� ���[�[h�LὍ�E`xД��ȢN]I}�vū�/�+ǲ�<��Zty�!�s�(S\�Ӫ��B�6w�SjX��&/��)�R������7��������������hܴB��$r�@X�����8�i��B��6�h������w�G��ґm^^r���0Y����jX�k1ܗB��#���_���h�U<p~rv5��.kG�:`��ֶ���S�~M����x��%��#��\�"�C�܀Cq�s�,\7"�H0��h�Y��B����L�d���a�8[�|OIA��^;��;���PwV���p��qqxK�'�����,w�C��N# ��-��m>���n.��V���w����k�<_���;��צ��{4��5�g4�R��#����	ܟF̊�TPx���I��Ե� 0�R���!��b����U��3���XYڋ���sv8�@u�읍�+ ��j�z�5���:��V?i��_�^�oV�:tݱ�`ZR*W?�߇�?{�^�י�S��M�d�4���I��<$,��C8,N��A�2�$;�U����d.;W'���X�Q�i8E7��5��l��<8�R�#z¶6ǯ�6�8���m��&��s�.��Y^D��,0=�C��nL�F�����s���㝈U�u=�-Uq׸C�I��?U���F�/D=��2h�cثU}�	qt��VR� ����2\��/�*[7}�8��S-�6ƪ�R*�nD���ؔ�/}Zl���7�V=]�n�H+��Wq��}�|.�@��7����@O+{�ȵ"��@l��Bռ����$v"�y���]������c@�.����A �<�[y_<�u��.i9��^����r�0�w��q�'�d�NK���R�`�ʁ|��jju�Uio�h. <�J&:k=e�!�.������
����Y��s�l�;�=����B��D�W�K��={������]�Ĉ^�	�o��1 օK�nO�*²�:+	'��0>���Q�#~��G4�hE������b�t.r�{نu\{m��M'>�^�6�C�~0�8��M�/�C_�H8uI��~�.���R�v�W)�9'�	h_�`�)��ŉ7���#�V�k�%��T���O񿝔����Wn�T]���#�Vg���p�/	^�4(�̮>F8V��\��+��c�OEKF����;0s�Y�[�J��쌒�=�>b� "�;���ԫV6���M�{����my%_1Yw�wG�m��H=�Ax @����X���5qkA�jό�pV����L�k�t��G[~d�ǚ��RAй�k��y��O����5�;�����1�|������m�B�0ŵ��tam��p���˔�bK���U���S\�r�B�!	���A�˧X��D�D|/�r/�� c�@f;a���&b=@DR�)��Z��;��*�(������7S��Ñ>V���9:��p��R�)GE������jO�D����G�{z���%���Ǌ��s PC�X66O����{.�AGqoX;�5��'����c�sz:i7��#D8��p�S���dQ,y����[��Des�5�lE��Ưn�8ow��G��׿G�%Fd�@��Cnsș�/M����:@�&�3�k5�[͗/����\~�%�m��Y���t�/�쭛k�ʓ�����@k�y�Q��';�mJ�3��v}+��o��;ⱜ3���wcS���4�9�?�E��!�W��%��ф ���<�Hٵ�� ��3�9�򚿊5�z����?����
�B�Ç��txǳ�V���1����ch-G��[J�uJ�lF��z� �0�4g��[x�~E*#@�#-������o�����A�WR�"����CI�~�rUz���%	��D�Y�[�`l�M�$����Юt����YX������%�G=h8Nf��&��)�8c���]�m/7��S�vɻ흥������7Ye-���>�vmNjD^H��gr?�����t���I��b�����Tz�ݐ��&b�d����,���
�RkϷ�W@M5�
P���_ *QL���E�8����f����c%����~E�f���d�gT~tȌ7��w�}�Ïb�
 ��w7~_�k7ڏ��"��R#�zc}�"�ޣ�ݴ�n.�3�:�eL昔5�[��2;?QZ��<���w�sTbQ?����C�,vˌ�g�c���h����6n���Sdt�(�Y�{�Y�� rͿ�7�C �N
nc$)�W�Σ!�'��/�\@�����|���
��͊���P6H��%1u���l���엃#b�g�_}�L��i���'>�޷�	��l�����c�����2?^��������Y��Ǉ�0;�5��
.��K�r�;#<�V��ܫ�\JR����:�[�i�{�������'���_��	[�
K���!�Ya�z�U�JU�\,͍�k��ϝ�4/�-��Y �5��BqH5��8�`�C���L@�i��\m���h/fVN�CT���/D�fݸ�Zoݐbl�ꒃ ͗"͞[R>.7���5o��tK�v�	�z>�����\/� =H�z ��F�/�b��/&�s��嘁�=�A1��OC)`�}�-�U�+��H�>�k`?)���{o�M6�l�6E2Q��Ƅ�3�y��j������2����z	յ����)�p
���[;S1Pu4HO$�}���ژ��2���l	�1��] 9��KH�i/���"�'7�j����D����a��G���] �cZ�%��p��i��J��m�£ɘ�
r3�~�i���r��t��G��f�%��\#�sBE� :0���^7�S;3PeiC�Ϻb�ԲN�|q�,�J�E�3XրW��o�%��f���f(��:��M7ɳľ��m�٭�m�}�����@E_��A_��4�ϭ[�>ϡ�%	�]��q@�� �ܪ$�G��;d�%�e/r�X�OL�r�9t��)M�m�3p &� %O-o�Ɨ��q
.�442I�6l��wOR׻Ta�,B׫�5aRz�T������n�SRaNK� �\��I��Z���ۥI�^Xc�7��s��ؐ�'�N�v}���2�p����s�%���l�i�	�M-������z�O:3Ag�U<Q�,�>z`��x4?�|��U�žE{���K�&m�����CC�	�6�T�N��*x�-�̽l��8�� $6@���f��Ń4�=�(SHEf�c6nu���	Cr� g/���{Wz|���6��G7�zO�dWO
�o�Ю$�H<�H�s��O�����\Zט�j7H�\�f�t@�W�bL�1�3�X�u^4�{?ڛZ�VC5<[bQ �oK��)�&��.�8[�9!H�a	��e�S��oFX;�V�G�O���n^')@1��@�ڌ�3�5��y����?ל��S"�9�O_�{vM�VI-�4@JMz�r��fK��9n*�h!ܕH�� }�}ey���lK��$��" y�|�nVO�&y&9�?��,�A��t���6�v���z_>�VZ����v ��C��$4ӆ��9W]��0k6�4�F/鍋Y�et>cmd��\i��a�*61���x§�<hT��)�?�e���F���r3��i3%x���8��R/�I�$0}y;*^�WkF�aB��Ԥ
�(��Ⱥ�؜�
=�)�㣑��$y�]/���>Z�h���A������!X
#�5�%1����x�n�FO�x�$0����[{�VA���s�R_.�x-^.�Y�? �G/hM�����Q��u���x!ug�����$N�M��(�����"�B�Gv��RPQ��u[w��e��5������u���AvԿ|��r<��b��S�>��O����Ĺ6`4��>Q�ѩM73�g���/B@��,�>����q�fS�y��d���@���ܔ�q`/��֣?�Cg s����s]���JΩ��Zo\���]���vM�����3�iy����0Fv`V�	�V3�[�
;H�6�[����Еs��4M�85"z���D��1K+k������]��/��/���m�=%]��}�����2�ٳ9]Ƽg��A �k�*��#[D��0b}8���~�Km�b2O�>�T��g@W��W%��e��S7��!lw�>����~ܩY��k��f{ͿQK�OLM���/����E�S����Ξ�'�	*�8>���Yx�˛�3�(�8n�B{=�t��wџ���_[� �"�b��oK�_�������E�VA�׾{��	Y��˥�L��*p��D�ʮ�?�ӣ��Ӓ�\�E��0������2�ޢ(�rZ���k%ݟ��D��
��ň�s�,��3�K/ %�e��H��iA�,�U��ǌD�qr���+R��1����Xq���e���.;g��ʂ*����C����N-:����d���욃�wŏ}��LV�u?�&��c���E�<a��n*M����&�H�\�b�~)`si�׷qz&�|�7L�5�[�O�̐����q-~m�	xC���f��O�Ȕ�֞I.�y�@o�W�l�f�ܜ�ѥ�~R���k@<��8N#S��ƴt�ی��$��j�|������v��T��*æ��a���i��1=�ỉ�m��r��"�%xk�����t��گ=)	�v#���옴1�2�u�l��^�9l�r��&aM|�}�퐜�h�K,�8��z�7����*���Y�BC��{�x�XH���(e�4(�(��D�~��=��`� ��7p���;%-?�͈�\�g]7���?*�b㘸�[ H�&u�3`m�УܾUzYE�y3.9�*(Y{��ԥK��k� ����.u+GR�o�I���f	�zC�iy%��P Pͮ�D��'at�wO��Rq���7A]}6���׾;��b�0k�����֪5'3�oMN�;ԥfl��%���[��y�q���U�C��y�A�:|��ί��c���;�A�-&�Ad%%�o
�(FGDO��n�t�h�(�ܓE1��
Q�}�h���F��ƪ04��d�U�`�q [��ˮ��}�*� �e���E�7�j�^�Z����t�k��gZ�?v�e�EG̲��?9�P�"��Ӹ�ٓN�����I�-��?N�\\�� 	���}������x�ּqD��m0n'�L,H��ir*)Bq�������	��:��t�-��D̓�c���TdyX�gEF�9uAF�&��צ��F-��g�%8�2g�/(�wV.�Qt���g�7-����^ղ�lpA��"���I��r���H���gG���Z*��1�p��s�?�s@ت�����J����\
�ir䐇í���nꇅ�?P�t_o�a����ßzC��{��aR1��.�8�QU�[{i	���`_���Â��GG0O����P�j���"(\�T�R���/�ok���n�la�+�5 ��:`��F�l��>b^��r�/��'nB_od�$=�&�[���6�����$̧�e���=��#��z���b�i�'}`ې>�vm�Qn���'��"�5.��JF e�S�2�����ɒ�-���5_�|J�ˎ���*RHY�m�J����{�^~ y��~��b�=�2Bǧҥ�>i��ߠ�Z�3s阘�6���M�)gg�LAr��8	���6@�$�@�(ȗ��l fzu�"	-��H3�+N�J�%튁����l�iؤ����+hN+�}J�3*�;b|������L��� �o'5�W�6��Qg��9Q�]W{��G#����r�nL����z��h���~o��k����&��'���؍�KÇ4 ���>��u��QzC�Ƕ�b�� T:�h�R��m��.s�g屡[|�<�F�����뒮�����n,_�180JVj�zt#�s�0��;L��z�'�	@
g�x�rW����D���/�N��"�L��e�8i�8{�O�(|PJv��N��~����
�s�~ݍ�ZAE�ƿ�LE�i�^�#	��X��������X�x�g�Lh�sO���T���|��Vk5
�]XY�!��w�5������I%S�@8��NX�G�|��q���h���Am�1�B�����_�a`���R��\ߛBG�-\�7c�l��:��E�c�c�'�G����U����K|b�2����D{�[�ˤ���1{Tjj�/�W�g�6#r�����9=ge��zP���8����
�tZb4~��]]��=���Ĩ����O`����k���wq��k�,G��o�9�ʍ�6"��ƙ&�eKh�/ܙ�oq�&d��W��>�������v�v\4�@Z)��I��K����a*lu9��S��N���Z�z�We��|�TeP��a��\g���fRj[�=U	a�P�R�͡�!n���᫃	`����T���	Ȟ%����]��,�;�4��<\
!�1t��X�G��<��6����.^�ǉ$O0����H(�� ùg��_���+�P \M�ه|��-�V8��sUB8�$��I���ֵ��	��\/i-��G�]QE�K�X�E�����B
+)gk�i��� 犈�p�$P������"�ke��ց1S�-��&�/��bf������7�Z�� ,�.H�h^������ry�j=QG	k�:�ެ��o��z�esq���	�
rpS��~��)��ӛ���Pjj�1~������uАJ>�qH�;�����u=��
�����#��{��&Pf���G����+���Zȯ�����a�����l]�,�~F�����9a{	��K��6f�����u�]��2����=��]�����u+Zm �B��k�$�U[aF�DZ���O��������Q��bT`�Y�
�_ǩ���SK<�J}�-���A�p��Y(�H�$�����H�ˁ�FA	_	���<���n���d�{܇)�]�NV�b�b�7P>���(�IA��X)j�y�+z}�|K\/Фy��سm�-��l"O�r;w0
<��/�
d����*�����,B���Z�;Y��������\��f�D=7�q�OKv����L��N�Z'�����[N��i?�����X��Tp�[x�[���e�n���T�< ��VA�mO��б0����.��
1p���	cg�gDN�c�/5N=�û�sygg�l?@�0���<B%�:�}�ܼ�s��2�O���F�z�����<оo;��t��)��H[��R�wR�� �=Me�5��ow[�i�a"?����ם��*֫Y.������tp���gvJJb�Lz	����љj�t��h��!$aNUb�X���m��sEv�h���4*!�8~Thʉ��?�͆��h�l؆Z��毦�~ä��8����pa�T�a����w��'z:2��O+�>$�ZPbl$��Q�C�Ea��7킭��C�Hk�s�?hZ�Ҽ���>�J��ytr;�ja`���2P/��l�&i���2I>����)��ףh��Ι���Tq��FL�V���8	c��K��^�I)7��*�`�;@y񏁞.l3u�OFM�7]?����}n8���S\9ˑ`�D$� 4RJ@�ٝI�U�>N�ht#>����J���[Z|���<�<�W���0���ĪtE��!4@.�� �J�$�Hͧ���o�	j��m���a��M��
�=D�
��;IǱg�;BBۚLA�ȝ߄�E@A[vҰ���Ǳ�ynT*M@�x~'��8�>�M�]�Zɫ3Z�V��	\e���Җ��}r�d6I{�_�!����84�r�b���R��Mr?��S�\�R$H$|q��(�'7g ��je�9�"	�5�F��y��Vȴ�ܞ���S(�t��X+�$��t��IL�庺p�a��\��k�u?�;����eR]�U�z��Cv�����q���?O��X�����r��|'�x���2sKLZQ�j{���������׳�+p�v�i;zg(��t�V�1�ɮ%��c�[�z������x
�&�8����z?��C[ZE�;~��Ф��:|7����t�{N���@�ӫ6F��ҟ!��v�w��&Ko���F��A�q�n�"� 3��.��r%@M���d�oZ���Đ�CDX�q��"6�V��oͺ��*do��Y���Η��B\��N��BK<�}��&�_�
+���p�����E_���,�&�����,7�Ҕ���{yQ�œ����sd��YЦ�T: б�D����]�zL�;����s��;�L�@�br�dPA��f,Ң���f�������+x0>����f�0��Xۏ���(���	�����{�m���*�"u��nfՑ��:��v��{��v�PBj�i�Icl�m�j��y)�~TZ�5N��{9z%�X��ԧt�.F1b�)�In���!��'-x��N�~l��~�Օ�G��yFI�*�����3eM�f ��\���*�\NR�| �pWX����->�(_��+f!�s�]_E��ٱ-&�y�w����coh�E��������6@��m��_Ѵ�Xo�"�B=�>J��]@X���{�\��?UL��$��qڴ�=D�ZooZ=���H�G�a%DY����V�C�P�zDgяU�Հ����!^�GZ��e�!9)��
��a�zϡ;�e��!Z�.Õg��Q�drd�_���L	��D�h��7��h1钲'e>Ʌq^ZF��Gl4H�5�	~�����C;���`t���#�r�T���N���/N����m�b���J����RR/�"rzmT~��8A���:�9��{?�T���<�[�xsc)0�n|4�*�i�p�=$]4!N����=�V�Թ����BJ�-����94��Q'D��._�������gthr�봃����x��\U���"�i���͘B���
������թ�g5��SO|^;�F�{��\�	�''�S_x�/�������:���1���0�@���&�bF�$]��ޱBvj][���Џ}�gߎCQLJI��`a��s�e��xS�F�?:�-2�8�:���f��X�d����B���a�XӺ�>��ǦOzF��^봃�.xM)���~�����6�s|*�]uAaLU��j��Qn�<�tNK`Ӫ���4�y���N��FX�T��5�r���T��A`���"��ʤ�i��)��թ`(v� �A��i����O������o�Q��u@�kȻ)�я!�d��6Ĕdب�J6�o-�RB��>�廈IeSImF����YwV����hvrh���c�R#_6d����}�@��� Y�vс���6�RBӢhL����L�P��k��QK���M9g��6��y\�7|�٤4��T�yԲJ�G��t�ҵx`�em!R�:D�&"-,�K(9`,���Em�9)���2�����Y�׺΄(��l��ĉ���
�EN��pGx/w�t%��zc�Z�9$���.���Y���I������&��e�[ ��ѣR��c�\�hӟ��$p��{�پ�N��O%�=9���8x�w��1Ri�$:�"��f�A���-�]F���i��'���.8d]�u�/E�y�?��	͏J��T�j�����Z�c�At�@��u�Ґ/���f¬ơy.�1���_��K2k�_�O��O�ul�AZ"�}�m�ś��c�
(]��R�''�M3�z���\b������ )+Z��o�Su(j0{�B�V����+K��������]S���'�/(Sj3��*Xn�
�IE���67�O?]~vKY���ej�[k�ԃ6����:b�j{)�{}!�.n�奣w�p(a�9Ǡ��-0_5��ߜ|�L�^2��u�*�d2�`�b�y���y���y.U󻿺R1r�`�h��.=絆���i!��d���jt���"8v��N�:�M(v��<=l��ip�?G!��z�
�����ތ^I=�0����BB�Tu��y���/>�ӉW���]~�zB4�N�2`��*���5�k�.$+����}����zs�����~�H��,��o�d�	G�We�.�b���sD�U��g5:dTN9�TL����0�4��陉�j���z�YBU��t�u�������T|>�q4�ϋ�M�=|˗�h|�O�W�*K�&� u��ʋ�Aq8���YV���fS���m�ʹQ���U1������[\�CP#�����xlB)���w��/l]��</<����)�ߡل�����0.I��I,]�#��U�+}�k�ĝ��Mh���M�%(�Y=8���㡯����r�����%i���Q`o"��:�Ie��7�\8\}ׅI��!��</%�Q���D�����^K�;�r��|M�8I�* �d��C��Pn�8�aOSgk�R��Rh�"�����m�T����A'�+�n�~�6��ΐB�#z�x��f,��s�)��������`A$q�)("c�Gթ��0�$�~L��,_�g�j�p���o�ȽŴB��P��b�\!_VX����C�!��:�^�Ɣ�`ú�W��X�Ґ&��Du>рԈ2/��T�m�)�Dj��b4�Ms#F�
~���Q��(��hn���-
�K*�0u0WN�sNPo5��tEՠ]v�s�!��q���)��0���V�p`Dq�1W���i���8ea̴A��ɱ���G����똫B҇ �>Ǒ�=�b�~س��'�t�q�K����2b4��BsG!e�M&���1|�ǧ1bd�g����+�LAI�a,tN%�@�V�8�4����@f��?~��0�����F#�ێ��W��µ^2�b��B�@f|���K�|,Nk��-x��?-� '�)�o����Q�?���G�n�!q�	���],s(�v�B�c
���v�#+�{�<�m�⡧� <��ASƺWl*+wu#W�#�Ģ�� G��o��{k� �U6\|�~ܲ�f�)�Ed'i-�橼����s ԃ�53Pe��B��&�K�@�%��ra��M��9�9	�\�S�u�������)F8��-�u�H�b�S �xo`1�T��=d�ѥ9G$`9�.7�9�%!��p���?ה���O��=^�)�`k�;�-����g Li�k� -8P���ʱ%��N%��J���j��auΤ�v�ޚ>M���#�C��5��R|s��D��t��tm,��]�R�vKLJa4�cx�(���,�(c�d4т*~�@�ZW7*�1:�؂�O���i-9���Zn�nYC<���h����mO�d�b�q,��F���vTS��v �d'O�����i�O;9��K���[��-#�� �AgG��8>��4ٛج�θI�_:���8IBI�*F}ox���j�O�J���yd�?"5��'����SͲ��󆍐��f�5�/�|��SD앑žzڴ[�%X��s��Z���5?ʹ`��W8r,>j4��ٕ6�JyŸ�,;�J�<�9�n��瞷��"����/�c�m(#v�i��~�$aJEa�݆|����v��L�L��/_짂���/Z��f��D~A��)���Hsp�4�7�� _.��@���T5q��S�9k��Qݪ^2�7!���;�VG�V=HN���F󲡑��XyA�m�P���i�'!�����:C��Hd����7����Je�Zb�KM��s�ǧ�<�D[�+D��ؘE6D���ݫ�s@�9*������r�E�/lW�H��!Oq�k���=���k�v����Տ����P���r%���h���À�>��@%|=1�4����E�e8�C�;���؛@p�\��f�憛]p���|���1;�vV��G��F7��V��`��������H2,-�ւ��d����4s&�m�cU� ���ֈI�'(q���"mXk,!'v�'�x[�n֭@� ��X!3S���K�m{�6��J���bKH�,��r��s��6�䍇�G���`�a7/ �����K���}����K�A�a��Č"������L|Ӕ��Vu�酽�d�/G�>�S�$��Pi��I}�=:>Y}����	0Ի�H�x�� ����7��r��Gs�(�5���ȧSf
���ۚ��{�ޞh'�I1^a��s�J��J���]Y�T��)�V�h�R]c��2�w2�v�����C�'�I}��w<;F<8�t
'�K'घT�	ە��]Cp��/�[�2����"[3���k���omu�dۖ�i���p���76�X�e_��՘�K(�Ip��$7ɰ�)	&�y)����6���PK?>�W�]�mC����+�IG��tK{�}1�W�SQ�K�.R[,���$�#�!|�C����1ԚYP�{w=u���L'�<�3�)��'P�,��	��J��i�t8~�eC��L��F� _��m����O2E�����?���c�@��9�XH٦�l"5e=r1+sQ1`�n,
�{�H����T�q�v��1T�>�	���H^	^٧s�6b�H���G�8�3��EWf%ِ�r#����txVؑ>��?64H=�����U�N���������/��G�}�ݺ�^}�Z�p.���^1�1��4����.���N��FM�c��|�U����8�/�֠�����AY�4Lz0�8����wMھ�A	�"�Y�VI&�}B�=�����gd���@������V�N20��`�I�׏��G�ssm�4����O���)�=�\�oZ`�8��avE��2Rg�F�py�A1��:���P���[�]vl ���5��?��f`9@~KkWσ!j�﹄t�N��I��kRq�m�a�م�
 pxiK$G���~䫺��E'i��G>݉�9l��'��B���Z�89S�~����^��r����!Yj��v?�������7�f 2��R�}@���O�KmfM��rțK 	W�[A��v��X'���N6H���� m��@ڸ�L�j�7�׽dV5��?r-����e��2����L���	��u��0яz�-Z�@3*\������S`ԫ�ܒ�rzI��}��?�(��}` &U�~s	�^�\�e_�d��$ܜ��wJ���B�BN��iqQ��RИ%7�@�^�-i��5��N�<�����	���)�|�7\q�)eȀ>�a�n���V0�b:��x���X���/�g����N0m��(XS��Q�UcD�f��Ϧ�h��?!�CL���������׿�`�kK1�i��L��1��B"2@�.�Śn薩�R���F���?��@�.�$Ph�M'�~>[��j�V�N��~��q���M��y���Xw��5N'������{��H���Pp�gH"��ƉT��WJJ:نJ�:�翘Q6������W��'���א	SCjlGJ.�m�,�d0�Z|�/�k;?�:4�;?����O�"��uC!ަ�Kݮ�W�S�׊b��|��EC)��'[����oжX����k�ַB�V�yNci�^�_��OLF��Kۊ���K�(1_�	�����lM7�����k��OSr���ea-$f���᝵��-T�P�^"/=�A �C�z���i���QYQ�d6o	�������F) ��X�}`H����	W0�>Tk�)��
����M��u�M��]@ᩕV�$��$��ջw�"@�'�Vs���c�n~�G��)�Rz�_�a�{k<���_KXLq��Y�Ҥ�<��i�á��a��l�$��01����E��Ҏ]��G�Hv���e~f�r�;�{t0��&�E�o2��J�Ѱ����{I���9�׋��ONm��)6]S4�
�gʅ�;�W�� CFP�Q�%3�P<��v�m�$m��d��zͳ/5�f%�q�!��_�|W	���zF�ፙ_0חj�Ďƃ?;�%f���T��zbe:�/Kss����������u���IY�7���,���п3���%ϙ]DD�ލsa
���x�'��_����q����;�j�+����;[L�!���}�k���~�Lڄ㜈��N�l��Qc�%�]|X����6����**����s�3|/!!fsm��I����& ����4;h!=�T��Z�-㬇���fQ�ѭ���JL3SA$�[.[��@��*b?�3u���cj����d�R]�Ci�h�"FV�%���Vx(sμ{[&h���#��H�Uee|��*ܣ��nK\pz�E5pg�B��8�2Z�i�[
�D�
W����t8:"*�T��D�7lh; "��p����R��p���P㽀����xط�^	l	ȓa��`R+��[/�e8�(�\����8��l*8R��\t?�ψ}�s�Ʀ��	�|Q���%(�G(�E�]S^i��S�J�|�A�=,�p� �/�����G,�'n�^چ�6Z��OdT�e�x����XՃW~�-�-����k��q|9G:��'�_� vT�7�P3v��<Ӯ_�Sبp����^�6���"��:�h������]vs$�o��o����J�N�o1iG��B���]�H�086��F��t�m����:C��Ju�AI,��ߌ�1��0]S��첄���H\r,�7����+�&���B��F�7m��&e��蕄�����cX{KSm�/���G�Gm�آϢ���~;6�<�,E�&��*��-�	�J���Y]��Qm�V�8�l~Ҏ��D�I�y�� W�- $��,?fL�~VHָ����S��p7	��[�#��'u1�Y��u�J�>����QĒI�Η���u�*�����E�!��Ib�Cl��3o{}k�I��]3��\���7s�#d<�@j�a��=��ęP����-nU�ߙ2!l!w�����t]`�u�w6��0Ф�y"����ཙ��:_ �%��9wc�/ֈ�%ݨk��cj^D�v�y�0l2u�/.�B�}1����?[lJxH*��w�7�H������������	-�Z�Lӯ��j~�r~��G�Ю�������u���(�f�(8��b�7G��t6Dݑ;@�J��속�� 4�规dD�=�`�G9l'�q����*������n���i0����r*�6���0��C$��>e��o�� ��5	�RAn�p�PN8o�Z��>oF�?
���z�h80�h���@M���m�F3�<��r�v� Ϣ����J�-1(ӣM��Ȧ�N��+TƖ���񒗲�Т4�b�3&bt���Z		���K��N�,��J=���#�I�����_����}�j�<8!,�Z��!�7�pW��*�iC�1���{V�v��[g�����0T���k5CS����3��7(��0�Yx3b
�#�$/���m�AZgr��ɝ/�����_u7�m�D��*d��nz|���`��On�p�ۻ���z��8�)��r�[�$�I�
���T5�Ck]
���j(|_,5`���ǻ[� ��D�g��-v	�F���Ǝ����h��� ���
��4pT���B*�@#~�Aօq	��k^ccu����;�;��`k������ۅY*��X�@�V
ѻ���S���/�2�M��P#���D^ԄY�h慇��?�r�Y�x_�-.Z�@|l��#��nŖ�����#����N݇���:�ݓQ��M����^\��(��T�M,<2���a�{!\��dכj�=e$���"�xO�_z����.�i��c��q������[���ʃ�������Y�)�+y%8�����x�N�.�~�8vJ��\��N��3h�k!]�"�R��s���F˅��6#�.>��L��H��m�n��P�&�
��C�g� ��֋U/��@����V�Lo
,�r�i����"��7�N��)�������R�����p�\1��˔\�k������딾�����r�l��/��b�Y*�ɹ|VG�7�8߹��
��p�i���4����J ���ǔ�Λe���._��ׂ�h��{�v�bV�O��9%���Urf]Ǫ���4ؼ�%�U`P�4)�@���D���z����Ǒt�_�I܀ _k@wt'Z=L��/�My�6��g���r�"�A:ׯ��#��'n�TM�a3%x�$�Uu��.rtt�P<?b*Y~$.��!:ߗ�EJyā���`�����v# +Ί��D6�|����u���%4�'5�­�Ŧ@�a�7P������3�G�V/�8���z�D����xu.�$z�y
?�?����:�=���S���2���;g
����.�$����0@'�D�kM����͡��g�+�5��T�$y=�*��TH_jP
�
R�1N���ד�Aa�L,D"ٔ��J�sbt+��\5|��/��`m���L]�pC�^n�lPh��pG�!V�����o��7*�[�e����%�{�H$�h���}=�$_�+ż
��x�( iW���J}׵_ ,M0�`0Q�;�T0��7�1�߬����O�!R��JY4,>Ẋ���u֯�'f43h��Z���"e�T�$'F�YV
�o��k\|�"Ќ�>]�(khEnѳ�m�)p��_����3��Kh$���_����S���C�g�Y��86�2q��~G'[+`Y��h@���
��ڋT����7���x���9V'��A�0��3w=���֌N��I��'��%m�O"���1Is��Xn.�I�� @�\�î���䅫�o�Қ���㪮�vg�vW�3F�����K�/�h���	)�Ŀn=��Q�CL�?�P�%M(����eE}xs���A$Q��Z@K�0m@�-k@�����%}py�ѻ��Z�����8+�˫��쯒��|�qE�t��V������s�o�0Y����kĪ\�J�B��$�j0��	D�\���5�ل�7N$H���aD!Bh�;��fzn���oh��)a+�Cz��1~F�C��*�	C��˕ jū���+!�H�"��bv��'�
r��|u,2��*�+Ѣۮ�^oRBN�ӔWQź� ��|��=K���9	��H;�n&C�Np��o��p���l:&+;��_8FA��pL�B�n����H�SS`���-fy{!xxg�߯u�80I�Qfu�	�6Z6����q��d՘k�[��8��׽�$~eѽ�M�� �R��@�ݘ��zٶ-ȯ�}�;B��D�ᄐ�tR��YՐ�uM?��<�r��EUa~�p���_y9�7�Z�$֮q}��hcv#�A��Ntt��{�M	���]��I�-tj�[����T'���k�Q\s�J���[Hkui=�@�5�l�7r�'^�⤷	H&b�p�O��2U�}���ߖ��h,(�&C�z�{r$��aˎ��"�#�3��c��l ,���c�n������p�&6+t�NDN}fQ�M���iA�O4�f��þF4��
�>���P�;��Ȩ��qX�.��#.�q�D.QKw���M��Uk��g9u�ǞM�����t��oZ���"��B䯇}�Σ҃#%�"�)����d?\��W���F�]3�G~���q|1���u���԰"LQ��D<y}����A�`�! ȥ���.~2��c�~P����FT��u����Ԩ��)�F�"��"e��.e�����d�8���m��a�����P�ʃ����:=�����}66�&�Y{��;Ӿ�!��l��8p��4Ј�vE"[#����-��4����'�w�t8��	�TL�5��p��_ōl�7�Z��h h��y;�`��^9� �|8�ܳђ�����+��e896�0U~3�V�<������{�r���qI���$f��ߛ��8jٵ����LL�#!��T�+��|Gl�y�e	�����(�3�G��C�����C)�H��� ���>\��B������hV�����D]�S��~��d��-�����i�K-+��a�����Y���y��:��X:jT?��_����Od���$�ly��x0#������ �4�x
���u�S@ӡݭG��Y��;������*?��� �:�q��*'�3=���r4-'r+��gi�_h��Y�[��9�A��զ�G=�߻�
/c�rE�K�h����	�	Z �Z�_�-u���-��*���|uD��G ��FŽa�J):��j������'��,uk`~Z�TW[<��Q@��}I�1^�^�~��"�.3��n�i�=�+��ʑ�����Y��S���/U�4���Đ~wz�k��{��N���+O�(� '��u���I�<IW��8SrQ��f�h��dBS�:5�WW��ε/o$_r��rч�oN��O�R���F9t�� 
�;Ȥ_�p�����:��$�#��h�s���W=�k���-Vc��� s�I	<�1��K�q�y�@���cG}��L�¹vg�sV�h��n�'FL��b�|ٟ|7����m�pT�tI�7�dk,�3���x3��U6+�h���FNo���
ݥ���_.�����*�6a��_��r}����S}K�%ƨ�ó�]�ߍG%99�Y�=7��S9a*H����'u2�y��M����[B��l��DM��S����Bf�0����)��ް������Vv�Dg7Q�	�a��ҋ>	�;#8�2�Չ�!���ߺ�T���y�	�	F(7=O��Yz��qy�(@���q���`��u_a����-#3@�v�ҘN���(�Rt��uǘ�-�W*��"�4A�<��^�(X�� �#CA1�^Z��y}�Dwo��5�KP?W�����W�������}�����9`��(R���C�[�N����?v�-�+��Յ��� -��}E��]�#������ҩ�gĦeF�ĵ���q�a{x6����޾Zp�/�|6[�wss_�h�SGW��!y^��sΤ���Ҳ�MB���e}�Q�D�q�{�A�>��
ҏa)e��g���Pe4 �t�2��4o�f�0���"�S6�T��`g��8F�	S�U���
�	u;��o���ܼ�M2PSAj/�|�ra<�تR��L>c����V�}h;�<N����-bHm~��w�Y���$����M .[��*�b=n*e��bwP<�;N3���)�nƷ��y�F�@���5��VD_����	��j��|�6������T��H���L����*/�&B��Xgɷd��$+�ծ衍���3���0��q���;;���D��j��#"M�as��uD�-�9��n���	N	H�eu���1v������}��j
}�ٖ5��)����6`�����R{�^ Te�U���X�ٷ�q��61��	P`CZ&Bg�Op3�郵o�����������:�E�fi_�A�~�N�i�4��Kj[�1+��W��n�>un2莑��lb}�ZM|�S�.��4o�@�dYJ&�.VPĂ�J�"� ����i�py��$��p�����NR�Prj<ܘ4�$aR0��&���/-b��V����s^��O�|��(�/qKt���%�ǟ��2�~\���m����a��x�u�՘05�������;���>��ѱ�[4��S�j��jq��(<�h-��
\�������]yr�x� _4TǦ��[N�Ph�߮"�N�LrF"�!�fS���>��n���BDjt��B����Iج�-:��_U)�`��ztr��<�KM�Q��D�����5=������3�h�\i�P�+�	uK�V��3C���~�����p�fӠ��zq�/G���:��d��y1������"��'�R`���m�&ig���9�Y�?6�vU!"]ɝ��)��/�b
�^�fpU
��ϧ����� r�Җ��b�7vĸǯ����^�=���.:�+P�1CN��75�����)��b\�
}�z
��&D&��0쀎r3Z	��D��#�
�BE����hf8`�}�R��P�����D�I�}��tR�R�gK�I���rwM�ɻc������f��q���4�Yv_�Z�WKf������d.�Ք�.l�ñe:6�P@��©~�n�·�nG�B�?���[c)�X#�󬰞pX��whv��#i�Xkr2���B����9}�,�+̶�Š�!g5���T׈x�|�>'U([XOm���KSG��*;WT�����L�MG���o�[2#�Ԏ�'cػ��N�����W�G-@�B���C�WS>��%�1A�8�pwP��DY]�5bXUm������q�k`g�3��tXLau�eg�׭�e|D�� v����Cm'���c�L��I}y,���@�އUq��Ȑ����
��K���S����!�Ag�
Q���8�T�؈�s�7N{�[�7�� [�ВF3Ԟ��OMs�ԭ,��!��D/Ɏ��[�hW:���çF2�^Y�d"c�2���C`�W�l6��j�Dej|Ar��1����=rg.�-:�ă��?����œ[�CSE��W�;����Ĳ�iP%�p���>�4
:,�]+
dH�"@��0oj�?��A��(��/zfa�"�s�"�G勬J�U_?M�����Xϗeo���/m���tAo��t�vf|� 8"�i���瘗xU���f��!��&�5�y�q�S{��/�����#��}�SF�#�~���O��\�}�v����O;�g�sY��#�� 0n�O�^���|�2n]�Z�c�u�eX�nZF��i�n�C$\$��Ɣ3a�����&p��ȴ��� �r\|��|��8���U��G)9h%��3�Tz�����rՆO�!B��\v15��4yu�����������6�5~��p���8_�f��� Zb��z��a�� �q�/���Bi�If9�28���8`ȭ���ј�ى� N���'��������n��M_^]|D|b܂q�b>R�����)�\��7Ε�_�v�.��)OU��h������}4�O#M8�	|/�;�˧���n�^�r��0�Z�=� žv_�9j����1�W�8�H ㉛Jݧ?4>����r�`ʓA��C0՘�[r&p`p�y���vׇ�;זw���d�}���}ݺ�G! 2��g�.��M�1��ll����;d�8.�h�Q� ����a��[V	>N-a���Y�ن�s� ^�u�=Yf�(�j�X`k\�Z������A�U�ʟ�)�)��6���D�|6P��v�|V�K�!.��y9��a���j~	��X~�շ���$Б���g�F��f��ƅ���1k&RN��A����*F���3J��8��$k6̢�c���D�׮�[�"gr��s��L�Q|S����1ʒ���ޤ��H�����D��ǻ/�4�;����)��|)�E��`�Y�AT�ӑ:�i.dh*�`ҋ����Ե�T�q��#/�Y�%2Q��zb��?��ޛ��7�V"M����ǿu.�{�Ʈ��39ՃG ʙz�ߕ�0�/s�>Z��H��$���/u�`y�w�y2dM��"���H}�I�.ZJ�l�f�"<�Lv
'n�uٶ)O_l$� $2������v\9P��_:��hb	�&��>�r\Ő��_�_N��v @l���؜�����u±q_�(�T��~�3�Ɖ����05�~<�Y���#�Fnu��s����}S푋���G���6�}m�R*�O�{&j�,��[�D��%.G@2tL�p׆��)�k�A�;��Ë7$KK� ������pԟ���9u֏L����0=��w���Ч���J�����1��7�eR�#Ci�$�i��[��ʕ{CuR<<vX�����в}����P�s
�^A�T)U�C��fo��JA�Հ*:�� ��;���%.d#X�6�)����P�}�����9+��h��:4ᙍr�.�&`��Tai�̤>՗��%�)r�G�/*����� ��JSqRO�D �)3C�J�Ҭ�g�E`f��U�V%?�[\�UE��9%�,OɅ�j���nχP��䝼bPf=l5^fY)�\�*P���L����@�\Ք��������$�(:[٣���ҟ��g��.�xB�~�6*��t��hqN���*�>g��=)$5�j̙y�'�R<�P9�l�Q�E��ޚ��6G���\6	��䤠�̶�xo�CcjF`�֝���ł�-���&*��p�]���	A�t�[�	?;Dd|J���^:<K���b�(��C�{��>�0I��;�kp��5lV��p�����Pp7��s�~>xȎ��^�L3B*���[���pi�-j��Pɒ=�V� ����k#O:*����.�L�D-t�cE��x���B�Rn�ۧI5�M�+
�Tbb/�>O�G���6�D+�"rZ�N��o�_2e�� ���AX������o�����>0Exq����t�_\�sV��a�#��=0Q�bd�\��*dn�����c�<H'g���^����o@@5���'��'J�n7F.��M��¡^�;�ZƔ<���#鷢�:]�@b��yI5�3��&!����@)Ԑ�+w5���2��d����{�^k�1��A�[�M-zgg+8�r�Y���y��u�Ay�Ǟ�����:1���rA� xX��fI����7�ɗ��.d($���{���H����L%�.>�:�o'`���&��i�������J��Z`�k�-66�,-���t�I0f���\��ԏ��h
X�o�!��鯑G3�u�hX�e?C���@��W��6�HQ^�g�xd���M+i��éI���冭�ӑ-|�U��u�x#?��1�$�+���lt�^	�eN]�_3�D�ʪiDk|L��xq��aT�o�6���9���G�p=�>=e�j/�ei���C2���SB�A���8��;��M�f�}�s�[�wW��{���4�S���[녟�}s��׮8�� �����C�-��L�܍�u�dQ.���m���u��x/�JQH��'��yA��s�Xb�B,�t�.s��;������	}E�����b�;B�#쪘0�R$�!�i/�����<B�r���٠�0l�PBe��'�����6C�N8.��`�����ᦿ�P�M��f�p�M0�=��9�µ���~����> }��^g�ᚧ�#�4P��Aw���$����᧜fg�4��$-��Q�R��l=f���P��ѪEf����EB���գh.ڹ�$�j7:5K;"���Q1�i���B��Ic�^vė��%������F!��D|I�ղ����ᚅظ�2�Sj#���k��uU��F{�=����� �*gt�s �^1`������K�[:�1ʪ��ܥ,Cڒf[C�a�2�%���b�Z��]ݬ�"�jZP�gJa �����W���75غ7���|����+x~8Ӟ�`�[:��n�
=�_[q�k'ܕZ�ġ(����Kd,�	v�6g�
>�'L6�!s�����ө1W��ٚ}J�sR��K|3�ٽb� �ٝ��|P�:Y�5�ÖO�'�!�zz��h`��˳Z�lf!��>Ձ��7�6��KR#�����_\�	!�n��^	�2���O:��q��Ё�[:��ψ=F�Gʽ�sĢ7._kt�~�4�С�H�0�
6ټ��n]Q[)����y�j]0T�-5z@���7�£9�`ߦ�����!��o��C��6I�.T����N�-:Cb+�m+E*gd/n �H�p���Y�\
�p�~��~|: -�(����=�.=�r5��v���?����b5�v9�ܢ�]�䓀�sD�~�>VU����_.��{\�5�V'8a|�(��&�ǲ�HXl��`.���T��#Z�/��O�d]�w��Ϙc����⻲y=[��>���^��q@�O���{�[��A����1+=d߸�R��-{Bv���qN>U	L��O)�)�È�i�oy\���f�Z彾���-�N�p���67Ѻ?P��=�V��fe�|��\=�V��Y�γ�L6m#Z���+q�o�"Ó��$=Nɿ"��8�e.����0�	��ޒC�h��XǬ���ޖK�J�����Ţ��`�S�����&s��L޿o^\u���C�#ڢ�k��`�Ku��4�A������|����u~@@�D�o�R��W{c�l�ŝ�t|g��979�?��s���5@[	�>!�zŀ}s�� �3����PR/|�l���_�-4���7h�x<�]��Hn����@� Rh}�i�p��A;�	!dW�q�P�J�G�S�Y��#F�
d���������o�;�	�|�É�L��ѕ��Ѹ�Xr)h��5����P��O ���"B��T5||%����.6� Y*!{�긞-�>�]���d�\4!^����6u��._��4Q��z�L�ޫ �w,Zy�t ��C�# k�5$y,�%��HV�ŵ��Q�%�/B�Ƿhl2�R�fu���=�"91Ԏ'����,(9�U~�÷f�BҖ�x�mjky�hTU��~��o�aFS����0���ۼPM�]umR����ΞrU+ܴ17h侥�
kD7t��T�}���	~����zl��g8>����:�( �3ꯕ�$�׭y޼"��M��@�T����Kj}qx�;�^��V�� ���L��]��Q���e�Zm���t���)½?�:T!F������P׈W\֯Ŀ�``��}��T5&��h2s9����؀)}���uvZs<���L��p���<l��������(�[f� ��>ޛ�W�:TZeq����g��-%"�<,Ʀ�ж��L�d�p�߆0�M�^[���5��o���wVY�%�ut;�u��g���	�3]@o/"	.�Oq���ϐ
����1o��	���)��ȫ2t&�����x(bCS����B�ͨj����g'G|��^˗g���
�����/��;@>a<��d۰��_�p�A��Gq�=�UE�W{�o~��YM�Qm��\��4�~0&Elw�3�3�����̥���c��Ie�}�E
�m��<��ȽU/�h�d'� ��d�=��z���BD�C� ������'���+�m!1�c��ѧ�Ҷp!�Z?��ح�û�?Q:���u���}N�F�cu>J�g�[���H��~*E'���$��.+�0Q����U��s���5��l����1��f����@y0�`��M�@H0dR5��Z��h���N�_+/�'`6A�ބ�>Ls������k5q�I;NI�zO"P�B��w�*�	����όwÚ�h�]$l�����ߋ?w0)��ݡ(���!W���� �$%�������"��q��e��4ŵ9���}�^G�8Oyx����~�ːE�%��������m�j�z!�}�=κ�hȹ}����!ɧ��=�"�S�����^�8�폛�9-��~:{��4#r��)�h��	#�E��*�u|u4V��Ԕ.����./��Vo��OH�!+,m�, ~�K��d©=׌h���V�����l�<p�j�Ez�V�riHO�JZ��]< �&oG��Kk?�Ȱ������Ϸ�	ALvV�͌I�,<E��l�r�V�	/#b�0�vD1ț?��p�FVN`�K�rه �,��zJ�'~�'�VT&�%x�&��ۻ 	B�n�δ�b����j �����Y����Ґ*A,��ͦθE�'�Uc�J3��K	�%�v�AE4�V+�M��m�*19k��s��ԯN�s�JrN�������L������]�eD������!�{��p���<;���C1���Hh�� gUc�Øu�5���s3���mK7�~���G��~��8Ӵ��**����f�-Bϫ���燂G$@�CAp�Б�Ҏ1F�o3���x��̵T�"�މ�>:t�Ϣ�b>%�v� ��\�v~��M�Α6�C�@.�o2��aFf��yc�(AƳ� q����&�� ~-3F5�?����27|�lN$�PO�%`	�t*���i�`�l&�b߭�������i���P����q�f�љlj�α�������_�h��8&�Ñ�~Z�aʾ�A� Dc ]H�$j��,h�Hޒm���1�F�kU�;�A�v��}<|�a<�\XV��P�!�P�~�+���6�|��h=��j��Q��҄�c.W��I��$�ӡIPn[01h�Ҡ�Hy�� ����|Z��x,��R"$��}qcv �"<�-��cwD�����J�fO�ōE���� QwH�ub(�Y��t��z��r��;UIF}!�uJ�tx�0��0�N��Y(��{|gZ���O����;2�݊�`���1�C���۫B������ӹkԈ��vAIZ�R��-����G{kh���7ѷ�-�П��ٜw3�n�����O��S�,��ŧ$X��5�-��椦Hqi�]�Ճ��S�Oi�t �U�p}�}���%���T�)'��B@�ʲ(���iOM���eU���[35LĠ�YQ�߳t�p���F2V�B��c����D<�|U6폠��	���l��%�������~��	�����eƮq��e|�)��x�g �@v�c����:�Y��b��@�D��9�X&���I�_.���8�v���*����.��hĵ���Rg]�u��������vP�[�Y��9j�\p���# �Ը=�����drD�by����c�z�� ��&����x�n7!���`�ZK�ßo}x0�3S�n���g��b2%pU�+M�ؚ�2w���p���>Ӹ^&�'��'��өC{���1P$�� �B��$���Xki��_1��u^J~l���:/B¥�0��L�/���hOD^)Eh<���fZ�,���kypd6a�/���zQ8��Y��l��`����y��,��ɱbA#�+���v�Xڈ�ߩ�A����}<��
W5n���t^�!�f���!�Ӧ��}}
M��wx���"VR�LD�����g�r�DT�c��ژ�qg:m3���
+�16���,�4�m��C�;Q���?�-�����t�6n���vr�1�'}���:���Q����8"�&��z�-_B�ScIH�̪p�*���_�����!�UT0]�k���)�g�4�St���w��,½�=9	gH�P	�f�E���|ƤcP��uCC�i'm��c�gk��ˡ�I��]���p�"ya˿c�-[�^A�Ζ����,(��z��GZ]�د���V\و�(�e&���}1v�E5
��/^n����?eos��={zfH;d��2
~7�Ҿ���tj>�����iJ1KƼ*3���*ׯ��qrx6����U�"|�6���Eұ�&)#��;�2{kr�%#�4�FA�W\��VGv���z���o���6�_<�H��U�����{t�Ɣ+Vޥ9O��:NL��ȍ�t3���9��N_��_��vS�)̱�£/�iP�L2�Z��U��[�=6,l��԰G�!@ZmLJ�(�5�?�:ZQ���$-��E⯨������xm6����^�I@`¾�Ib��rKVfrOɧ�R��]R�ĆK0z� �]�H4���F�p�B�.��`��O�Ѷ�;2���;j���?��A�8=�tH�j���]��п��a��i�>(\�_Cy}0�uZ5d���s%.��_i<���2�l�.���J��.��{�㴣d���U��|3}4ư��J�[�(�*ڟd�W9b�9�O�X��	r��v�x��iv���ړc�Ec�"V�<��Hb��~���fK��c�K(����2佾��~��.؃�~�>�]��O=�qJ�^��J�����W���d���Xi&sg��V�2�	�uL��'���nZ����`�h��;߉*��<wN�H�q�</�O2��ѩ�/�d�Ė��7�a��
+�'���w�A%��W�%��K�u&vz��M$�9]�,�jEg�@w�ѐt�/"2_y��N	�v6�(ػ!�*pt���������r�-"�8�|�1L�ɂf1r�_��W�;h�V�ӯ_�{p��m"����c�e��2�ۿt(d��ջ��~��=���44t�M,��1
���б{�KmF����Y�<'|��G-yh�Td?���%���T-p��?9Z�z����^^��C�8y�c������|��.z�žr�����QH-������_r��"A3���[7t~�j��0*�J��:�� ��r�����)x�I'�C���snk���]"m�ܿ�t�r�/���g�_���Lg<A���WE�|�L�HW.�����]�����K�y���>�Y�"a���ztD�|�&o�����,	�L{h>[�G~.Z6�:�K���e�����D��(��nҨ��P�%�(sn�>�=zz��.Wswd%Eāc5��e˺E��ul�lbG�ok������f� k�3�������P�r ���^��Y���Т}��+���.�:��Fe�:w�!/�4�:�䖬���0�	&O�Ư��b't'r�ۍ�LB�%^}����=��4/����z���d�2�j�\��r�t{,ѕ�Q�6JN��^�W�+���0
v��)A��}))=lkguyF= t#��1��n�J��0���R�hF�H�=�'�D�<(�D)f3L�U+0���!��ק\���
'�u��������$�I��5�͎qh�;gs"�"��׍	j����w�����+G�,�/}ɾ(�X>�"ڐhݖ�F�2�R���u�>~������;��fx��f=(�u���ۉz��$'���P>K�Yj2=����:�d.>��_�윴�Ndzf�2�>��,s-�h'�a�S?�BRDfY�Ҟ9i�|F�$��ֶ�����V>�A�"Fy7�f%�}��`_������a�̅_r0졛�;�6���5�G�x��0�p8�n������&��0U�m1��.{�\�Ǚfg��r骢d������V	EZQYg�����W�4�i6��2�9	=�k��G���^���!-r��Agt=�J]�Rh�a�z�Y���Z���;��
6]�լ����:��江����	�N�M�rٌ��Q�:Έz�e��F��R�l,qI3~��[P��=7���T�OrM�D�_������m�1�ӂ���N�Q{R�[l�My`i��_7&��M�wt��t�������a&I�:�(�?�JF(��*���ہ�2^�Z
�#�EKƙ빌�fp�v
-�!�����Ʌ��=�sg�O��$��2��`�����Fu������e'��޼}��¼��<�;ZcM{�հ�m6? ��~����+�wt���Y>uVBp�H�t���A(�7�b��<b�qVk�M���t|�pz�VּȰ�Іgnx�z���%��k�U�
cs�bw���e�e`).�]{�
��Oa?��Įae����+����J.���j�����༟'b��p�tVl��A(�Ճ��ȧdLp�*�m���g�qM2���Q
z�K��Oޫ=&L(=����4���̠x��]��\0m�F�0���<βDQ�GFa��g/��_� �%�WX1n����V4/`�+|��L�6���x8��cv�Oi�1��a�!�{q%q�d�{Ħ����r�U�Έ���S($�&@`���h�;�`�c�vr1��j��j�u���C3�[���L��x�耝6����3@MH:���oid��-�^V~�bN!�����N�6Pƶ�?�M����3�.(~������m�-Qƃ�?�-�,聈e�.k&0O:_Þ`��y{&?��M��9�OŽ;*^n�Ďv��"���7(A_������S�8t��z�k��Щ����"�Dc�Qa��m����k���LF��6t��"
1�I��3���,�G@B�1��?~C^�B]ϛ��G��F�h�Gc=�� �8&
���
X(�-=\� ��`��=��K|��?+F�jM�K �@��9�I�p�b��#�m�v�"=<�?U)ʞ1�8DZʤ�י,�������u3��ܫV�15�l�Ƨk ��~���F�rb�fZ���d�����a���/�.�h%�Rb.�0=J����*�
x��`�����V��u?2lP������k��rb�m�2u)�����Q�(M���;��A�6��cd�[���$�T4��ex��=F����*;�bh�)�t�Qo�O'����rc��`�ⴷ��D�7@�����[F?��]���"�Bq��+�R����5�z>MP�{p.}���J]a������V�O$��q�Hj�����*��r��+��ʗ�q[��u�� ��]��\Â�+%�Q�Y�nW�vϜ��s��8fE��=S�	�8���!0�u�xI�Y�Ɏ�z����w? *�.����,��ph����'���ca����/ݖ�'����6l����(��(�U����3�S�7�t|��s����[BL������E����6�;�S�����j�F`XnH
�
��8�̟�(���a��CHE�q4`=��񔔦�< P����;Yr�{-g- v��e��#G}�.�	B����2�bW1�#���N�ym�#�{����q��~	�YՎgҖżD�#���m^�\sGHߟ�4���m8��ry"�F� �v�x�t\8S����C_k�I�Fm9�T~��o?�W�9��#���9�W�_\q*��58�_+�����X1:e�8wWn �U>�\����s]�A��uqܙ��r;�ܘ��6}�Ց��U�"9�ޢ��v��!d|�.D��Z ��ô�6	I��>�Y /�-���EV_$L{����n��8/oz�������u���*QL�tY�u�N��La"@���׫�j� sfDn��1|� ݮ�n#�^'�P�P���+a,��H�����8���d��!|��qA��	z�f��D{��gV(��xp׏�9^=�����B�(o��:���y�)k^�}=����m_	d�=��lVص	;7yu�.���ك�����-ia�]���*Ą�P�p�� B��5�7�,a5.����u�3�D�?�I$;?����(E]3��t�N]V�D����n&�3eɐkم^Q��t��\�4`ħ/,_�q��?�9��w��e��LU�cZ_&F��?G�aPQ��D�1�A����7�Y��QK`(���4=�O�<@W����zט��Ep=C��o�]3��]J0=,K���G��������0wm������F,p"��^~��5D�_�w�g���0�VcN��'o+OM��l�,�x�Ʋ��T�J����-�:�c�B!S��_�倗	�*/��ýlϦ���N[0Q�i��h&��Ŀ���j̔�6sL(����jn{U�	8C����|@��W��r=���Or0������eS���[Y����WD�[S�x��|��)�E�Q���������("\uC;��g�O:g�H~VG��K�R2n3�v�%�f�L��}`�3��_�D��RVV�g@H����w ZŧS�(>R.n�=c�v=oV��Z��ާ����D&7���`Tg4��H�TU��4-�Ӆ�|�}2*,걮wJu�����C 9"�v�g�4����P�\���!�_}f�G��������m���|`Np�O�o�?�;�0;/�(�qA٠��� �(�����4�{0A۰�����dt0k��he${�v&�}7�v��`�c����Ҽ����œ�&U�H�� OREv�c�'���&FqB6S�R�����lV���ZѲ z֟�v��8�G�����d���?�D���*���)cx��Ň���_JV��$�cJ��yd��'����J���&����c�$���ec�kI!<���@3��6���M��:�t'?�/��t�#�h����
)w��'d�\?�jt�{^���,.>��&���%k'
�@ߤ�|�]�ټjgŊ�E��n5bOz�Xe��)k�����k2ipBz��!���C��_@l�v�yn��A(����<��b���Ӑ9Ȗ�{ۣ���%ڕZr��I�&[���,�7��P�gq�+O��]�RM`�B_t�5����_!m�&j��c$�4n��<�������[�(�'��d�^��0R6O���mUA���DA�(8o)���0��#+���|�ja3��-�"+)ט!�S���Z�	s��"lV�my�ڌ3����ɶhe[u΄N��0��1Q$����(�ڳ褄���~�i�.z�s�8�ﻭ�
�s���kX�H��l�Y�
!\�x��b� I#�k%Pӓ-�2��� X�^��J��7V�5
���XT�z��],�Oք�&X1	/�Z;\gC���lc�9�P��Ғ�5+�t�5�9�O��T�|�%\G�gVe�;i
z�%iѬ�1�K-���A�Ê�u���v��je�x�4��3�h�w�pZ��Iu�j/ r��+�PT���]�I���~IܺT���oN��r�yYf}��NRfl�y�uc�h����������%\@�H���q"�otkË��Q�d�l��IH��x��C������;Ֆ�b�y��S�ex��D,i�A �SW�$��>�V\�\E@É�����g2���(�^ad�s]!��lI�,g���	�~p>�j+wE����kw4���_:�VfJ+e�p]H���`�)����	�Y��`EJ���|����8�U=��q���Q��y�9�_eE�����\���a���i�	�G���ܚ*�#�8)�x�\GӨu�d]?Ą�&�]���_�FI�/Лy��_�RNV�A�4l��j'<�Y�H�s��N%l+�F�>�Wt�M�?ńa�B[*qTʥ������-�`�V:S�u훻7��G��T�`�� �,�z�Ba��0�i�>E�h�(������q�o�H�J8<�4-�wR�s��Kt���UtE�!�$�)��������Y/��<���x�3�0��.�ܔ���!�Ӫ�2��6��G��Y��K���hʼ�HG���%
��G�C�8;Wn
nb#
�۞p �4� L�4�NB�K��Ɍ�?���������������2+�o�W=�u��V��'<�1�1b�T_P+�㾒��8 ��l�-+�<�6��x�4�M��c��{� 51�W"$��tg�O�ͧ�*�7Fȣn�GY�W��`9�V�������هr�I�5+�5�T�z��&�V��S⳥�d��/�9���T��Tׁ|8�����
T��C�<�zCN��,Tc�&���m�N��ђ��-k"'�׳tS����A�F�K��H����K�|8I�4� f�������h��������YKv��,|9�x�3��x�� ���Ԫ�^���9K�*5�g��^dS��ƽ�z�x&d�"k��Q|r�P�l^yڧV����:�5�e�_=��dS|�ᄬ3�,:�MEX���r@�)�Uz;�$�,�? �� =$h��i�B̗�J�T29��:���U|i���T�@	5a !�%�`�'���󳵲#� (����h,�ō��j~�����v�jm�4�2s ��h�Z��]���y�8����ELP�/��ω��0�5�P�c�/ [kle�a���vx����˥HC��+,�]b��_ c�.n8�I�Io���+���3��v���qF$q�"O��U��[�21ڡ�E��N��
W�4)T�bH��1�q��#��t��;$@yq��)ٜ(�:���e�O��}I;�+�]�Y�6Y�?,�:�3NoWޚ��d�2�9��^H.5'q�~O�sի�Y�����G�1ڶ4�P�����sTLNQY��aUf{6z��TI=Wz|��u�:^�n�3�XN�\B^�rW����:�EM�NV�q��5*���Qu�e�oY�������x�U�ʆ������N����W�l�i,�l�����rou��1乭S����p�*ldP�\q�R�����go����/�^�,� J�������+驩��u�W�-���d$�E��U�r"��A��P�ӲD/uqG�6��@6�NY���3��<d㸵�F3A �v����F��P>�)QR��K�\/��B��;Z2~X�_�҄T��D��g�ҕ�x �/N(�k0�h����#����'���AK@�������2�C�����W�9�OKf��v%+�� m�S��vƤ��}ԭ�Z�"�6���.[r�
�D!/ ���`lJ�DZ/�EL�{�QO��7��7f�q݀"�J��T8o{�3w6���+�'�i'{�ς�$b�9l�^���V� �yB�II�b�K:	tǉa8R�]��!�+���;��}II�����N� s�H����/P��(��󨣸~�Z,#3D	�����A��a/��/�3��.~q`��8�ԛ�Ov�����'1f��ќ[U	ˣk������&W���ojN	˻I����r<�S4t4��L@%/0v�6v�
L`�NHb��k��7�A�v�r�8���t��t�Ē[+�)J.D�P���&�\9j��qd�o�n�����4���F�(�F@�j�A�)c-�C2��է��`���m�J�e����*�Sp�TA��#am�f��Ʈ���ܦW����4�zS�tOt<�i'JsΎ����	�P�
C�`���8/�8� �_�>��u�&.��,"<7[i���L˦�ڴ���,![jjH�u�|%!�]���h�f~�]>�A���@�<]F�1b��+y�)��e���?)�?�N&L&�X�f�)u�θ��}���O�\�-gy��F(y��s���η��З�nD>���c��*�)���>�"���˘���<!J��)/�o�ks�"8@!7bl���Kފ�(2�܀���$��d~"��2��R���6���YE�Xo�6Y�����Sc�?w�Yy�^�ہz�	��j�;m��2.K���E�&�9�e=Rj��&G'X�	2�tbu�kH�X4쌗a��~�"�f��i����+��s����P8N���y�	T]5�A�ی9�4�a��|�v*�n},1dң����}Y*>b��O#�鏪vZ������
�7Hk�)o�d!���*�;��d��O�9������ڱY�h�����sۚI�Oj=��=�ϖ.=6g�!u�K =R�00<v��b0C|�c@��{`����������<�*Dw����aM1������dud�	_�����w��;���
1��O4�uF�B_C�u������[S�[mMG�_�Xo=��!��6�:�����\�+K���+�֜xKfi�Y�IA�y�̡�����e���sF���`f�#ՙ���s��������4`ט���K�^N��y��A$�aE�"�&84���HwZ!i���NTm�1��]D�:r@�)��Qc�L@��k��d�������3��ӏ�Co�$��9rɍ ��Fs�l��;�h�:Av9�F�@a�P�$هذ��D� �l����t����y������0�}�{n�P1����@"�������{`t���jr�G;��*<*��L2l�a`�^|:���k�oT�T��ibW�@�7�����	��"�ӻ���[����B�����L^{Z�r@G�9����@���e��͑�:l����g^���g��+�Px��Ը�w:g�貼��x�?�%�PhUXI�@��L3�;Z��q:C�>�$$���E#wJ+��"a6����2���H�o:�E�{֜�Zv��t�'=�3��̣���m�)bQ�l	�G�Ha�8ۏ����V���k�ۥ柎����M+��tW��tq�R�d-��:�K܈8����H�U�zK���n��2�ip�̷��qn��6�,���bU�x�x�9C��t���F����.d����z�B�n�-�2Wdun���153#9���S��P�׋ܭk�s�g�����x��\�YB�jE���>��E�|��ۥN�(d�I<~�.����16��6-�i�,݊Z?<*>Xnn1����R����Lgv�����(�����ߦ�i�{Qء y��~xC3l���s�/�8�j�񁮤W�emI�̤�H�f@O'���z�6�ͦk*�P�d�#	<���|��p_ZL��XR�?M���� ���oL����X�Z���G�Iґ[hh�w��qv��yw��0�σT��b��}/��٧�	��]Oyv�~� �UF\R˞�v�%�}vF�#O}س�{s-{Xr8��X
C(ī�f����.��BX=I���:xs�8R�7�FFC5Ma�6���__�����JU/~�܄Yq�'H���^��Z;A}돦i�}�^�Z�=�ьby<5�W�râc�3�y(H\gd��+���a��=E���+P�p\�A��w��aQ<z��F*���w0Y�����K���#ڢr�j�W��� 0��ĎY���d�)���b�tk*uFh��p	#��'��o꿝���������bCL��	�V;δU��~Mb��X��f�(Z�9v���.���j�*\\�2@b���c�E'���2�%��9�8�/����ڋ�q��@�;딱<���w{�X���������%زr�<1���ᴾ��힜��ϱ�u��uv��2|F܍��z����=8����4�u=�~1f�'��ߥ��a��Ph��bi�� �7Yq`C-p�xG`�2���tw��|�@�#z�ŀ���]�A�؂	��T��;�6
g��m�����1��|������s�].$�
|�l��H��il�>A&��$m���_R(,�D�g�������Ta��Y���D���m�i�� ��P?��nn�M�FzL��� �Ы�f2d�{ƃ�u�0�Zr�z�ѓ�������[g��e�;s���rn�_�L� ��`����iBS`O����ϭpK��2���#���	ۦsx:�.Cl�nl�o-�2͗:@��������/R��Y~�'_���o����XJ-���6�$�4P��T�N��=��aS*ø�E�H�g�-z�\�P�@���w��|?`+]x�:v�]�a2�)@�yJ��xF��������[-��4l���R��S>��^P�(%@st'��j�"v�R�u��y��&wx̹U��%f�_�J�C��[)t�N��veit[�k�t�K�ٮD[߫�oS��]^U1,Q^�ov�gd��!ɫ��l�ẜ��S>,{���/� �ދ�N����|�҉���bL�TF݇j�
��`U�8m��ozuB��L�=i�
�\ �<<OKcG�j1��<�������dI*��l�T��>K�-ų H�i�+�i5���p#��q�����G��I��c�JI��B ��%�:��4mA�S ���H"t
~�)U�P�{˘�lB����ƾ���w�q�a?���6{��_ɱ�-�U!"�C
���V�h�'�/�(8��%^���J\i�򅟊�<g��M��S��{p본�+���r�U�I�EV_�����A|��B=�x`V�د��]^�k�_�*S�����֠D��:X(%�{�U�)�)D���
�k��/�İ�*13e4��j��衪�K�q�>�rO�N�G�z1�2�r.����+�Z�e�r�݆1���s��9اȀ�`��}�O��D޺#��3=@��A��k"�Sc�����IF��y����^wi����l���?�?���͑m�N��>�u�`7	�Q*5z3��ŋ,���_6"F�=Cy��d�G� �ל�m��Iz�m����D�/�o�i���QI ����ڥo����[o�q�l�g���Y�����pV�j��"PMHH���߼��Ӵn��ܽ��qV�袏ROc��Ӽj���"d�]Q�xt�^�h b%������k;XE��3�^�������>R��+!�%nYl���H@i!�b�?Uz�E�ێ%ʈ�H��H�g�4g�d���N�0e�����V�/U�a^;��G�4,@�Dx������B���o��A� ߣ���$7��>����)l;��n�a��l�����j��r��� ��Z�-�[���$�(T�517�R^���Mnd�'~˾뎩Dx��N���6|.C#P�'T��I�F��ǚ����f�bɿ�T1�6Q#an�8�Q�,#Ik����mRk�]���Nt:� ���WH�5��7���e&��Y,6�R�
�E�&"�u�˛,Fʪ됡�@��~�fЃ�K�*�أ��`Pid��O�J��<lQ��곍هH꛱���3�[9��¡���:��m~Ko%�[Ճ�ihx�,Y)��@X��Z��W�ި���Vp�o	c�!Lak�q�L����`S�ص�;����̵+�r�d�Ƶ�f��[�a��ꮁd����m��'����H�_�:�Չ�&C�;;dY��{��"7���hä-���@I�&� y�Zn�ث�HR(���j��������O>�ķ�N�R�W��d������,ݫX
���Ħc?������mA,�X��ܲ��:��_���lm:���3�N��0��:��׫4���)�y�:?@+�P��ŷcx��1�[W>���#� ��T���S�?\�zU�3�z֥!�d�9SEؚ>����GT�Z3�S�	hGN���`�����4^ >�����[#��+ }�;�֩����f�l���
M$��Ҽ8M��늏�kW�ayrufI����X�`�έV]D�Ȏ>[e��^�2��S�=�{^z'���O�u~��
Z#�ٕ=�z�?�ʼ\�j����4���ԛ^m����r���`
*��ߢ}E?3����c/�6H���`n�+������ �S�۝h[f�[9pQHT�S3�.�����1����rJ�F�Aܨ�:�4ؤ����;@:yW��oh�ڥ���u�,p����a�wНB3�6���$�E��cw~&�N9^9�S�����Lj��WT�.wG/�������Ad8m�P�sJ�"  �a�u`Z ���D��+��n0�8��c���|I�gP)��iSձ�V��؂pIm4�%|�V�1�O:@c�	�]�w��nE��h�n���ln_6�Ơw�&�0����Z7�A�D���n>a�������r��ge�2pB�0�V	f�Ep����P����c��T��c����'���{HY�^b�f�"���?О�t����p��b1K���tׂh�I�M�0w����+�($�ۥ�,��������/��nW�.�\::�t���,���$��%��Q�1�B[�S��@�H�d�muV���"JH%�����s��t0��O�ee��C$��f�'���.o��N�=����+�ĠJx�ת�� (Y��s�q�}�7T��\� �*�� ��;[�I�ٗ��S�?�⬢-�@_�,��)
_�=����z�f��G,w}�}�89�ǆ?/�cw�V�e\�y�}N�X��hflV�!��e}k�R�h��e�Vu��`|嗘��0�nvE��p�(B����\ph^|���O�w]}~A7"-�R���_9-�����B�f�U� �����c���\�
�B[��1� rw�[H�:�K;�z�2�cP|)p��&q���M���ԞRj:E?�'��@I.S��x	�
{��<���������㗺ّp���J�Z�i#�W$P�EuL�f�s>���{��E}�c	[����o��,�N��q֧{�����=o��t�ЋJ�ƞ��U����,a;,2�}����t�XkXD���H�FY��(z��H;y(}2��z�abT=oq�Ȑ���=�x�y �����U䰢��+o�~Cf;�"*� 6x3zH��f|0��
vJ谉}z�ۋ���ם��
����L����Q��bDXf9��;����i�!��z���f\����N�D�}o5g�5a��e�X�=z���[�*`���ʫF�u������&=#��ױ�mK�\�����)'&�X}i�vU��g�p��i#�/���]�M@�E��
᩵Zğ�C>^��%p�mN�Z�L��=��e�%K�"�r�k���7�c���5?�}���C���2�2>�=z��z�[f? ��)�tX�?�4Mn>��X?�ϗn=AW���k�L�7�����!�dȌ@��lCF�����+C�/�娪-���0�9O�%y9�|��덵ɡK�>f�4�{o�QƓHSw1�t����D����k���k����y��Ժ���0^#m�^as��z.��!+�;ɳ0+��(����z"X]�(-̏&U���״^�_d��C�����t�\���#��&�\��L�,��R0P�lϊц���vk��r�Z=a��3k?	�5߶b#��a	\S�٫n�X�U{6����a����ۅ�d,�7��,$y�o9o���-��	¤I�����k�*V�Һ�u#Y� Ǐ�ٹ�%�V���`ADQ��|��4-uO���Pz���?��"�4� 3ʸԸB��׾/�D�� ����Z
���-*~.��klem��Ӽ�Џ��6$J������}SXU�����8���;�����[ǑeNSK�X6��7�sGK*�LF`^=!P��c�v5�U�Wӫ�ڠ��w���P�H��rk��xK|�K��b�Y�s��c����Kf�T3����씫.[�5�߂�ޔٝ�[��߱��&1����
�H��y��$ü��PM�rQ'����>���/������}G�qn��HtQ'��V⥾n�0d�L7QfϤ�s�����Q+��^	��la�$}6ٜ�B*�����A>G����]�g�Q	 �y�ڸ�lZz,�Z�������ڒe���3�_Lt��V�M�z�\���J+_�9�Px�.�r#�F��� �dӫ��'�4�u覺0r�%����]����E�e%?
mɬUc�7Ͼ���U.	,pͬ9�v�7��:(@�|O�`ZdyW�!7��!?6)�?d��o-s!?�����E)��ɞ�8��Q����4��1 ���x��L���5�آ*�����Q#(+!<�: ��c	���Ƣ���_MTc��.�r����:#Y�8U.��Bt���}��E�z������|�>:we3����R�y���WK��/1�`��[V��-q�P+n�u�pw��0�A��(�h�B�;�'�=�L���լ����s�@��s�6q����+hk�	������(��pF�w��*_Վ$��?�m�E�ml���"Ø.�]˖]람�����w�(}��sL�_���EW�b��ت�w�t�����.��ĚΫ^�`і^y��Ḍ����.����:h�Tb?��D���;=5h*6����baĞ�R*�9����
$���8"�z?�1�ҶV��������r<_"�)SMU[�QQDL�����ӂ�0g+���1�$��u\�gWi�M�s��.�qoi�~��·#q )��� ��%�ɮ�."z����<�Ϣ0����UI���&��P�7-�ھEp�BmP32F�+xG��%N�y\��p��˕藽&#b�ʌ��ߘGg�բ϶#�PߵP���GJ0�@z�%IAdN�K�$�V�@�WR�o�(U+FX^����@�s���&���LțM�*��`�q��"�p�/���y��()tu�th�Q��^{���mYE�����8b����!��e�w">��18�4+0�z�]�	�O��	�����^��i�8��@�g��Fo�	���
��/�g�/��)���Ai�~���śX戦�,�"YlMǑ�R��]!���%�F�
F^�x����[�q�G�9��=�@�8���o(�b&u���F�r�����*	S��>�e�枎(��8�ų�m��֐�K� >m�wO���+n���� �F�;�+���{��vŵƃA���k���\P�@�m� ���X�y*�U�b��|�`M���ov��r*����۝z|I�	Ȇ�+Vl~�<v:�
��%����)�%֥�4�C�?���%c�:7�c�H����0�Z b���e,�٤F�S�E(���~ �-��;��w��0�gL�f�G�<�lPngЁ�ɟ�g��9��nj��^-v|�n�v�����
�	7M3P��w`�<��r�2�2�|@�[���5��=)J����H�C2F�>F���?VJe�6���F�ǻ.mv�k�΢nU�v�`�И1X����8�Q���pV�;9%H,g�_��wލU�O���f�Hs����[�&'���fJgrU��8�昲�k���d�����|g�SS���M=�Ӥ��I ���}���-7��}ڟ�s�I��urg~����̆v�д�����4�����G%�~)> ��:;�K-Q�D�*jN�@�h������,��4.w��?@�A�)u�N�2�w�?}������FV�	��u�_{ݘ�!��n2��.s�6�ԟT��WJݱ׳d�	�nPR�8+�O^ڎ�I'����:�؝�w*t�����2u��8�l^N��.�=z*�� �i��_�E�*"\�Kf2�He�|Ե/����]Q����J���Z��Ѳ.����p��Q�?��m�1���W�Mv��ߑ�1!V7��H����� 6E��5 0���y�
�ŧ���u7I��bɧ�,&���w?���
���6�AE�^��ttr�p.�B�46}ȭ;<�#�㑷��k�1 �N�O��p~�u�}���VCg�����a�~��	�A�e4�U�B���\:�NRtY+ƙ�/�bےbK��DN���n3��͵�y�����fV�H
��
���%���C�%5�#���1^ppͷ
�ňt*�<*I�6L>�)�H{ 8�寧��y$��� �c������7�(���3�7�AD���[a�w��?k���
�����zQ�l>)�֞G|.���dB�1���0�]4w��7�ٛ��� ޢC�һpu&���}M$�?$h���x=j�ɒ�h��jI�b1��v�zt��}��z�ru������	����� �S�9A9��M �$t�T��������	Lk�q���}Q��@��!�9,+j�f�g�쾦C�Np����.��!0s���^}n�xI�G������ ܸ�6Bmس ��iqnWRخ@�J��0�r���BYk����[͙O����2���ܺc��*���k)����p�E�U>`��u
����PqoǊ��y�:y�>�A���(��m	@S��.����?W	<|��MqZ+�N<ȣ��-�rRy�B�0^� � �߹U�
�?��"�`�D�}��$���U���Nj��ԤM޹��|�L���m�K��JI�{��9fMn���&�P[B�32�R��7Mq��E���I���P�g�/y@a����A�P;5��t%4if��R��&Ի*�	���djO��	2U����Q��K׃f7��oB���ˍ��B��(@e}+{�!����w��t�Ӵ�U\�1�G����`�k �7�HL3�����#�|I�ts|�j�h�=e#G�l�m�f��t��*�k[O:��Q�Ӳ�O�1�3�9�gixgy��'g���O��[V�7���u򞖁�oxZ¢�.���`L�����bΑ����k�����۾�	hL.��Py��j�{^��A+�U Q��E L�"��M��"�L����Q*¦K���{���������)���1ޑa�>!�%�X9`�)z�5���H�����G��x
���D$3T@������f��\t�����W��W��d������3�j��&��2(�ݪT��O��Rʰ�z=�Ks������/���$� �V@��\�6'Jl��A
��	 ��!ضao�i�Ȝ�K�p�Z�6�p#�F]v��d=aj(�ۗ���бiEҾ�r|@�-V:]1J��l�������tJ�ƋR�&��M�	ê�^*oI��5�A��ͦ�i��������6h8;���4����rr�Ra}�h>���To�Fc$+�vT�%��7	f$_�C�Ye��Mk���T����c'"Y�u�
Ol���r{|Ɲ�s�:�4�M��#�T��:f������zA��!�k�Z�\�v��6��l��-�idk=�Ā}���'y5�_t��)��K�P&&9�>���U��y�&UyI�fB��b����o"K�y+��=*чF�����Q����Lˢ. �M�n+Js�������I6ݷ�.��h����7��ꧨ�S����ߒ(5َ�[ɠ�W3��#
��z�8$��Hv�]�*��U�L�h���W��q��G?�5rޭϿ�p��u�t�1���d.=���%�E
v|Q�)ůQἾ�VS�N��}���".��hm6T� 9�$zf��_�x���nIo���H�p�,�%9��e��Ģ0��׹�ˎs����i֥������!w��,���H�*T��^�!�|��@����z�W�٩]�`�
���x+����C�7�x��Wx�&����c�J�.�U:��V�`SĜԜR{��A|aUq� ���n x���]m�i ���Pލ:D���0A�6�2���P�R!�^��BA#E�&�I��9�et��#+��HE����;��'l2�WLE8��N�i6���$U�}/O�.7�4J���5�3�q4��W_�PT��p؃o�0E�r�����w��B\� �{@��4������7���^<>c�o���s�o�_l*�ρlv���d����}��o�_�kg�o�n#=��['s.���,�9St�G� Y���B�q�����6����W��k�֨QE�Gv�$�U�̺�����蘌RVk��Vؙ��>O��/���J!�o���E0���5�ŝe0����yͪ���$�G9�i�+$"1�B�x|���[p��6���ꤪ�,�ҏ�jX���Rv-�pE��!OU��������u�6dh��}(��;����I��&���}�;�
<�]������-q���ܯl�`ԑ@�9GZ�=����9�屡�U�W_f]��hk���/��:�������?g���@��7 �~	+z-m,R'���\��ݚw�5	mﰹ�cx:������� k�������xY�-��0�V�T-u��s&U_a��~|�u�ɱ	Ƶ�cJPd~fe),Nx��V��emO`[��V:�{�j,�����wd!la���r�Ao�t�a��c�����g��j��Mnf��ɹŧ1��z�j-�#���$zEYCA�{�ۧp�ś��Ӡ����2XK��Km�}�n/cw�I 8!R!�Me,���c��m?��;�_1�l�Ua[_Oe�c�{cCƮ�к)�QPz�r�A/��	�Gݐ��T@I�l1�z�iQEYYn9OH�Ƿ�Ä[�K��a��?
!��pA���1P%���Λ!gr�,���'�ͦ�H$4 �����.|�{Z�ֻzH'c�er��V���Mo��R��8�r]�^g�Mix g��ӹ��aO
!
6L~DD�`�Qq����=���0����
�9ӫnr���cM����s����ʏ;����4!+�p�#�,��[�Tx8�!�T��C�^������(�Q&�9��0)���ϗW;�&v��D-[.���.���C��_�ڿ�I�a`W�+u�F�%�j���KF��7*2�.���ڻ$���Dj�΁����h2�gN�p�ӄ��"Uԃ�e�ٛ�����`O�[�K!������̌|~�l�������*�R��{n�orט*M��,u�~B��\�g�Z����=�G޶�?m����U�μV���֫�Q��T��)W���-,T�:^|݂�4�KKV%�5�2�?�[4	���_��� �NY77\.gm(���*4KN�kɃ��;�������n�Y^��ko:�I�j5�"�5>��<Qo��+d��2��k��~�/�J��4V��j���+%9Ic�ͳ���rי��V��׃Vc�����g'<u��?w$����� �l�tSP��<�_���4#P��0�8�NtK�&dIL��W�2�/1j��ł��(rċ�0c�;�'Zl��Ȧ��`��g�H��ҙy}A�w�o	S���x�+��y8�&&:	����c<C���a�s��9�f ˕B� 'Lǁ%� �Lk�A����$��[n�{�����@���uK�<���ruL_�8�oKr��%C���9��������[��̕�n9��
����
2�f��p`�rz��#�<�y�B2!��ݴ\vooA��$�R���t&у�y
�Ϙ�	A��b�[������֩�LPb�ʡ��M�`�y݈�)Ԥ_�_�ZJ T�~.�$UD�(�z��nW��$˂G�:e4ף���d?�mr˸֋��@e��R���^�)�x2��	�y�,/hC���H;�4��srF��T��A������_�$&SCbTy��V��F"w�m�*��`��hU��;�I%��f����׳��y��i�Qi �\ka�F�����vOa݁�Ԩpwp��o�)*���E(ul���ZN�M}���H���Y\���Q���ġ^<t��/���;Y��[>ZS��oBH$ҽ����7���&�E#�|���K�+�&|�+���#��l�S�!�V�Ҡr��8W�� ӏϣ8��:��8f�@�g����H�%wK����Y��@p�tْ4����J+ب��@C砉���j��I׷5k⽒0Q�y+{S�s�7'=(}��-�%��yV�^���{�;k�ݺD�$Bm)��n)@&%�/5hʤ5������,͟	0"#\,����k����[����*���>�j9hp�X{dIK	V�+/���V��xj@��-�ڱ�q�v�����-�+e����
Ǟ��d> $��S�y,��M��"��xO)(��(	.�^�J�o�f�-wi��p{!Bm���Y�Bn;�� g���?
������v@-�#����1M�ﹷ���7�j�ݽK�����±B��g��q��;��*@�g�J����?�y�k ����
��#�B��_��vi�rq�+"e^��tTY2EN�P[��$�z/I���Ȋ��K4���xb�g�@\����q��Sa423C�����F;&9;<��P�j}��@���7�{�͠L�j._�S�ULHɬE���0�T��d\3��
�z֖���^�Eڐ>[@-[���<�t9�]S<��pyjX��q�X��N���8l���Կ�~���e��=2-����J9���"���*�zot�!Y�ZR��4*��KX�Ek�}�x�}���� ���0���U���K���j,�ׅ��d%��/=��7݂�M*���F+8-ϻ��uH�Mː%r�V�IFW�I�0#�������Nͱ��	��qe:T	��=kh�u{=R�F�!�Քl�SQT�#{��M�Rj���{�io�+�$���e�U	ս�p[v,~ Rrs�G��X�}�?-{q�de���
�-h���{��Ӭ2��j��䊉`���l�jJ�.%7��'���"w��2{^�^$G��� ]�[�\]���hK+L�`y�����A�*�u��K��Њ٥ͅ���@2-��F�d�I��!���풴�|�ǣ!�W>����Bֺ�+�q�Q�e�_����G�	Y��=�W=J�Ņ���ϰ{}�/kdk�?�K��⑛�C#��j��E聧^����y`q��>Jp-�ǅ���-"��B��}��i%��X?�n��� ��v ؒ�a9���@�XV��$i|)x��/�4��&^iA-LD���`��I�{´ǖIp�J�[�@�ɰ:f��Le����H"ǰ�QO8�2=t`3����I"3�Q(o�G��*�p��Tn�����كaO3o�R��V�]XV�k����ҨN��D��Vy���m�tE5������ �<�Ӷ�RZO�"^�h��_�I4Jp��ȝ�W�bv��~��y�ڰ�N��fOז"�4Iy�T&~(@voQ�D"�(���5��Fn��*����vP#��Kx�&)�i���X"�^A��9Pt�`�N:�E���+�3�χ���n��Ǥb3T8�_���+�E�&E�̝3�����P��a���=x��BM���=;'��G�ǵ�P,S ��D4z�c/n���Χ�J���H�\H��R�E$&�0ﰓn���yk0��	�
��Nb�YQ�#��X��Y�4AO��b]��n9/�|���x����9�*��޴������B�]��B{�ʾy(T���W1d��������1���Ԟ�cm��iJo��a��yx�	4�
I�����, �c���m���]}��Jq�:E~��M������1�c|�i�W��YdC�T�͎vJa�e�NQ�R%�SeU���W]�u-h1
�x�{.�,pD5����İ����_FȖ8�g�3��cG�hl��^sD۲r
�t:�>����ޥ	׳ÿ��>�ץ�V�H���8<Ck��׼�������v� �?p9�[��{>Ŭs���'`�I���pH�rP���h�R����&?:i��@���R,i�"����?��v��b�K+�ޅ��r�Gξ�m� o�Pe���<{��h�X�&V���d���W��A�&��bZ�ڬ�l���r%�Zҿ�Ɇ�@�BN	(9��-hز��r�Jg��})}2(l�\4��G��K�/rT��cK�WW�?+�����5YJ�J�U�uG�����;�*�fCdeACJ��sc��ؘ�g �c��f	]�
������Jd��"U�=4V�s��|,�\�Zj9�FA��-Wf���]�ɲ]lR��}����b���'�|u3h��,�X�9³2B�0Hf��NB_\���d͂�qZt�CE�K��i�˭�ѻQ^r�����Ջ�g@�5-E�#�j��h��>�1���B��8r�2���b�r�iZ;����t1�p��޵�{Z8ɮv�d��8(yYe)�,��QB�˲W�61E��HrZ��Z	�&��®⩱=M�U���S]�W�'(�d��ot��C���]M|����t��@0�?미����[�垅�Y�_G�~�>����_�R� 0�_�|%a Z���� [#ݴ�z���=���͞�Q�)�JHF,�R�<M�,����",<���,�'���L�om'�<Q�`ܺ1Al�a���qӲМ�` �Z���hb��$�Y���T��Qh��T ���zR2�Qb�����ɇB���k�R	/�,^����Bo��N�y� P!9�}kZ�fý�b��>�g�1<���,��uY X���hr"3����� �]�b����ƚ�to��Z���d�mڤ�r��1A^���"T�Y���r���s/��Q�@˂�~��m���Ò~8n��_����VL���տ�D&���֍��Yz�#xt��7x"�rÙ�Mt@j���\
��*�O���e\N��'�#0�]��u�������5��d�5?��c���W��e�[i�T*�/�%��qn*XO|귬0���6�0^j�+l���=q9�!��
@��@�8�H�6�ߨ�Xp�8�r}�%�kv��r�����^��YꬮԢ�|���EO�
��D�E�����sT�k�$��P��g�� Jsx�����z��?z��k���V[����$�_�-���9�A�=j��ţ;b��jD5M�h��}Ɗ:n]f)���8���ۄDA&mV��d���m�5Q�wW[��>wV�h�Q?�Z���\�����t�"�x��=��Z@z��Yz��H��RR�w��[s�t]���BE�T���W��{��`�3��*([ɰ��k:�)�_%��rbS��n���q ���	�;/�/$J��B���Y0]��]��%� ?�H8ۆz�X�Aٯ~����+ �LD@c�BT��a?t;x��L�T�����Ɔ���OmV�d�Zt�����ν=��_aD��|�-��@��Ͼ������7=J/ě�Z������H�N>C����i�v�E�	�=Z1��w�h��5���=��nӔ��yF���b|�Z�k���w@S�F�ZD~�ixO���֣�2xW:���kb�C�矄��h"䌓I3�I͗����tS��P�� z��Igf 6���4��ό�p�d�i�(���QFEK�W�����eK��0K
� P�~e�̻hL�����Ӌ�9�^��!�܎^dt�37ܲ�2q.�ּVAC���A�b�"S�j�B����,���V�C��>r�n��:��0܈Y��?nI���ĳ��B�ڷ.Z������R���Ք�
7�W%{��C�`M���{+G�u꣩�6�U�Qag"���.��&%՚��T���y�-�cG.��T���{�Lz�!1^�C���mH�f{��s��Kn�y�l���2�S�st�s�� !)�����|����	(O�K��/>��QM]�`Cs�qT큢�f�\�8�ڂ��S�[ ���rN�"�|;�Qk�FA��w���eL�HUn�(o����V�I�0�R"�C�+�#C���R��O�Ƕ�'���BL@8M�~sӪ�x��Z���ٚO!���$�:?�UQ�z���������+G�Ev�*���O�<sC�z�h��%ҍ�k/m��V+'g�)�Ra����
���f~� �ttO�gu�/4��/C<�2����ṋTb��(,���-EO��E�%���0�a%i(��?莔b�f?W(�5�? I��H$��cAT��}d�k��3��+��=����	;�,^m �V��\�}�cp9���Cyu8���J��¥h*&�y���俙m�>�X�w��U��GSi1?�s�[��Á7���nO��ً�[�\�q�K���P����r���W��dn�ƙ��gT�R�;c�"���$B�����M\�H��W�De�śQ�<�Z����c��a�������ډ b��J��D�vµ�&`���px��x�����ل�t�鎾�s@����/H��ҁEgo!V�O���4&��Y>�1�	�P����&����m�f&����[l�ܳ�I�)�0�{2���w��1�c�L�lP�X��Q��@
78�G;~�`o��� :�t���Ԟ�1�����o�Ԙ5'�~#*��k�pӿꄏb"~	oT �i-�� �o�5l��C��-L����u���S�|��㷌@�6�
IzH��܂�%�[���>7�Z~o�m�������Z�N�
���H���&P	���/b�C��]�/�R-�:���^բ%3D4<�x��W?h�@��s~��P�-��A�;��C�
�p2a�7* �����"2�Ï%ӕq1�5�B�e=��&8�.�u��u�V?͊0�H�oTY�9��4���j��aH�T�H�� ,���E	�<~���0�3�UM�� mht���X=h�y}b0V����@���t�'����q���>���a�ay`�T��{��o��s��k�C���z��v8(%[��o��])/?�Cx��_#Uw���t4�BR�5#�+(���y�Q�� GB�������%��X�X'��U�V�8C�oJ�񞁫��I*	����N��@#��ݿ�B�xd�_-��%j©��=��ᙜ�E��.�u���g������m�X8:�J~t���,��0KUA���Q�G(��?�s��(�����u.8`���8M;G�fS]3�ke?b1��)���� e�W
��\��9ѐ�e��d,�N�B4V [��ȸ���Eu$Z�k�l�]ԅ�;����$r�A-�D�����eJG7>�q�p�U�Va��e\��e�fn�ie�՝J��ܔ������ĠZ; 6����95sVC�p";q��� ^��Y��R]~^
p�MAOw��p�\�L����&tڽ�3��3렻�?_�j/��I�������Ȉ�G�fu��
_� 86�dQQG]�'#z	�t 3����ɪ���J���(;� c�3��S�P`Z6&��.�f����s�CF��'H_U��|��/q�����b �\��mJBi�y�w��nz	�bl�:,��5G"ܶ��T,����J���^r��s�-��/[�
��~�V�8�_�g,�{'쁝�{N:)���z�����2���9�P�}#��T�52���	JX��6o�1��h���ՙ_���v���6ɸ��՗�X)���}7�u��"+�HO@��\s)&rʈ$�tƘ���ލ�������~
�/�~�S��h�HgP��lC'H�E�V����&0�״ �]<���ܵsE�s�K'�K���'�S�I`,���׋"�J�D5�2���@���j�ɳ�So����PB���IQ��[)Dע!�u�p����9rh����d毢+V�(���o�n�T�����3�V}CC�<�'�p�⤽��9߳�Ѐ������š6?h�}��=6�An[�_��ѭ��*C O�����_N��;�G��K7�Ma�*�P��B��Ia�7j�Oc{z$L�ѕ4��'>��
J|2��"�|�׶Λ>	�<� ��(���G��Ja1}qB�����(}+�S�,��T��k�w�I_��E`�9!'����cqX���3_� �������4/׊&^|R]�z�}�M���\S$/w c��kp��p��]f�2�r��ŭI���sX�p�MD�Cl�Ћ�5~Y���k��Di�AFP�t	���fNȝ�67�i$4�'j1.Fz���lL��u��@�0翗}S��	�͝Y�BSK�.a��9qF�nn��G�)x�`-FmǴ��>d�Z�`G������8D`"%e�\�J����K����V���&@D!�
*�����v�n�tmẌ́=��hw��}B��X$���WO4��.�y��|K�t�P��p�!�ך�a�=�j����� �O�.�ݦ�e�U'�d��_.I�3�����5����V��IA�K��h$���@"w�:_b�p�HC����䋊�	ٍ]���P��cf��u�.��>&ƀ�����տ���G��kR �<�aD��:��?�K3/8_k~�!���pj�d�*Q�����������_@����ʰ_�$�z�R�!���X�� B_�-+��
Ugc����[<D\*�K���i`�men�4�3HӮ�l��>�L�]�9Q�	�HRÝ�E���)��hGe�tq�ʼ)�żd�����Ш����? �L�ٵ��oσ�2Bu0n*<1KK�AK����ӫ�"�[�C/7( �K�5�
�+2Z즞,t�Z=8qXF̘-{8�wo����)v�y}l�4q}�A���%�;�L�Gh�|�#�Ϯ����Z@��3U���@l�x	�}���e�]��Jj^���f9Zx|Ѿ9�����i��)��6ٵ�	W^6ݧD��!ý����b�ӳ��]�΂����y�T��v��A��ih;a.es���o}���L��^g]�YP+CB�z�Ƨ@*m����[�[Ԏc�ϝ��Pf�A�e�n#�ճ(e^ڢ��i�c͔���"Z����h�f���^�}C'�>ר�Z�Oɒ�8h����~'
E
wZLÉS�9�m`�QQ�:��*(�r4���ߦ�q�#����83
�_��o���p�@i#X
.�Q���jf	}�~����l^��_���{S=z�E҃yk��Q	DX�N���z�L�}*��t�k�y�GT��$��L@� %�|�d3eҩ�p�x@����XTA��e�� =CaK޾�t� �hf��0(�Gx�ޠ���]�_�-Ɛ7GoN6����E ��0��5���f͆�Y�N
��0���R��̅Y���Q��&��lz/����w�q��gOH��R~�["�O#�@�9��ax�bD5�f�S5�Z�Tp�E�%w,�690��q\9�y�i/�� ���ҡv���R��_ ���⣏�'L�԰#MY���z�ls&?���M"��^��r	�Ǜ�)�:�
��QgEW��qEדN)�Mw�G�����'O{1;�@���̷�[��t�^�f�bPӗ�t��v'z�L<Kc��o����k,��3c���I�}���f�3��&r��[[z����Jz��q�zWEv޾4H�-͠�6��8�͈{y;Zʝ�C2��3�i���0.OS��S�;�K�M�5��p��.��e�_E�=�� �O#���� �c@�o��YN�f���u����_�ow|�����anc�̯.uK!H�ۍ�N�w�NZ3Q˴������ڃPL���Y]�ݥ�Á�YJ�{��i'��g{b�d.�K���*��WW�Y�؛#����pu`Z1l\w��	��I��(��=�6�i�Ӣ=Vn�u2��ϳm�,.1Qc���x�؈O�W�m�;�b�IE �np	�{���W-Q��&a�Ӈ.�m}�*r
��:Y ����U��j�b������[ੈ�/oV����@h�ܐ�B�-U��f{��aȲ���К��	2-�{v�����[/)�6�'��ڵ&}�Gk^��XDN�x�a�@�JT�*�r����m�N��Z��f��G؏�]�W~g����	�J���i8�.(�?U�!u�������Y*���������~OM��j�(�)������A/���(qY:�G��V��P�ԭV�YÎs%W���n�v�	n��VZ�ڥ�5`ի�TM5����8���`�Q��9��zw���Mi����!��:H�M�4~.��;O�4#��+j�9���HM���&�j~�饹/�����z#�tta��w�h\-���$s|��nP
>W��@��#��[$)�x#�d:�#���:
X"l�a���F*q���Z����Ӝ!)С�\�U!�̵i��K�3��,�A�f�}/@�";�	��,���C)��H͢*�y�WT�J"��OI-|a<N�N��p������4�`�G�|�u������x�5,"%!z���GW����'[@�E����}NfX��8Ώ���mf�i�'6�ڡ�Y\1��O$�=�Bڀ���SE���I6��}�$�-�� �,CQbE�a������3���`V�q�]J�����˪W=�l%�Y�0⸃u��\����8gIb��Y���8����S(��ј�j�(�x�����/N�v�O�)B���o<�0�qp	liƄ�^���NO"�]`�� ���5�}�*zdY�J-���>����p��}��>iqH��O�v{A�m��OY׽�S�m�#�8=|�U��酪�J$X<7 [
���Qܦp��2ɇ��;b{L�횎��~)0�/���.ה	yHf^3T�v�0�p��5�ϘiĨI��j k��K�f~��R����L__��u���μn���I�1��(@w���g��Ha�QR�_���ÿCu���a��O�K@���nQ�^���,�b���㳲|�3ri�������@�Gg�1�Xj��:Z4@]k�Y�sM1�nD��0F��(?$d�T��Iې�-L6y翴=���G�p1�F9��,j�8�ۀxtDU�h��&�}ce~���=`V+��%��r�FKv�����x4
�R���ť�J��5:�-�����F�&��*Yx�~0&�(ϣ�Ĉ�
������=�����?��I�-��c��@��OݺWN� u�4�\��Nv�G1��C�1�����e�#Fگ���G��',{;`�Sd4P��	|k�������Y�鏵����)���!��駘�_��Q1�c$F���w�����&�F��@�tp��f'�Q�C����]�B�w2z
!e�'�WH��_4OO��#d��K��-k�`o�)4�F��"��Ypi���
��旸:[����b*�+œ$�>p`�)��x�Z�Om���ޮ{�Ɗ^�p�z�]�~R}5���~�`��!�N�%�dKM�؂R�a�G̅�r���}�½�}2��_�ۨ��v= ]4�v8w�����>/�Uc�v%���L8oQ}�lx|x\*�v[������hn�AbJ
J�m��fÕQ�H2��K
�!�1�܍���k=�+��fO�r��T�݃QD�vz�r�#�����ur��yС���,��`��:����7y�%�&S���0#sU[%Ԫ-���!���~�%ʁlf  {;�0�N��? JL��އ��u�+�qp��_��^�5�L>6t��z)l_��=��j2����I�OjD��;�k��J���Q�S��JF�]�� �����Z{z�]+�(ڇKW91l^5@�JռS�R���cr��Q��w�di�Фd��1���2���;�KD)��*Nz�N��x�?�����K=-�ᛝJ�x&= z�ք��^��r�y�;�4MH��K�qjs��l�t�pt���[5<����r�w����svP�G�_
@�c|�nGb��nC9���������#��B_���y�|3P^�x�.	�G��ԋ0���,�k9-��'P��fU3��rx�wv3�/�gXE����@ʬ�(���ѯ6w�C?x@��8 ��_�\�Q��12vBM�j��cݠ���F��oɁ�`�[Jy�Q�)���?
Ơ}���;M5,(I��'���KB�98s��Y�m��n1��ݑ��D��׻A�����|�U	-9�Q��l��<q<A��43~Pi7�i:�HsW}��h ˭pUL�@��u~ �3��O�Ǆ���,3���Y2@�}���0{�b ����?^�{ }��*0��B��B��
���K[�b�)ˢ����0�N���5���,��烔u�a���Ľ;�-�K?]p��s���3���5z�vJ����m^0ر��v� �~Ě]�!D'ݺ�$��޽�x\�Ɓ�I62�ОÏ*(�˖��xvoB��2�^�X���ٳl�9Gc'!��_1��B��.$" �7%�0x�u�d��(�5g�2��~ŭ�z�.vә�Hy'=���쩼Q�4��yX8�T��N���1?�w�ߏ���_UW�'�2j����h������Eju�=�A��_ƙ�>��yzZ^���'�I��P��D�_րz�H7�z�m���ɺ�M_���fr.t��xzhI�f��>��5ȿ�8�vN��^���M�Ke3�%�Iﯗ��6��2oح�if|�1\.�_�O�_2yS��u�ˍ�����r8lX�&�1:��1��D�.gCL�Pӥ��q+%y���S؁x���Lׅ=��l�s �D���t�o��S��|a���g����R*��+_�C��6�C'�ܐǷ��$ڱ$N��>���M�_�3�p��I-ZM���R�fx�f��1�^���Y��
̃Ƶ)rjW������|��VnY�E��������a�-�Zv�idu����¢��������'QJ�|4	���ЭQY��V�����^[�-�7�L<���ܢ?�@�>��A&�;�����)����s0@,��Lz������i&��Sf�-��i3��Ňx�c-6"�۽� �q�rÂU�6@�]s����{�L��ȬԸ�wOm)�ˋ���!B�Ì�U(�M7�[m&#����z�e�ԧ�d1~�8Y
;���������a;�����
M���*$��h�9OU��'0�eh�޶p4c_	�O�{������ǧ�����TvH�_�@Qg:�!MBc]+Q�l�əE����5nPԔ��#F�+��m�U�2�d"�4�#�p�����	PWj>Ó�Z"6+E2v����Eu'�2�j�C�9�f���m`ڳ.��Q���^�?݄m_(:�p=�b���D��� ɝd[w8��ݡ��'K�Q��r�t��i�3����tZ����B����M�2.�w�meB�Y����>����〢�oE:4'�I�t�v�Q��/�혈e@�O^aVk�F���Dp�k	���C�.+/�P�$!/��9���ŷs���K�	��U������Yk��-�q��v��J0��s��0�Q~�n";��.)�B����j��+�K�Ӳ2�\���-�w�X�n��,�e5�񄌫I��H�J Y�b�(8Yea"��L��р\J��-v�4���c������O(�B��C�������O� ��S 6D�*.�Ѳ�YHR���'��E�I��=]�>��)c׊t"�}Y�[����0��ؘ�.�N����߷�ȇ��dL�'z��">����9U�0፹$�ÖR'�2?j�]<�14pVSy��S�5{����o��+����.y���=[�󻾷6�pj��2��0�q�9��gX;[Ds�?@��U<qk(�Ʈ�Z�@�:N�F�����P>�R�3��?�!�vn�)nS������ۂ�,��8���1b�u7b1���Ig�w봡�m[�,v�S|!4�9$���=�����jhx�Y�]�T��󎵙�-���o�%+,��D<m=>��kq<'�o(�th�;lzb�8��J7������k^6��wi�����cS��+�
@j�ovlĴ������2N��F#R訖2�t�mӐ��{"J�؜z�{B�|M	.-�8�m㏃	d���%���І��A�+m>Q�t��F/���Մ��o])�#[����2�N �g�z_�9�g=��ӹ�O�����iϔ|1�O��Ǹ�?v�.Ƶ�+2���ь01�#.��\�4�#���=n�Y7r��S-%��n%6Њ��K��S +�;8G~�X.�O���Z�-i�B��?�װ�FcUJ�@7�S�T{�*�f���s��P�3J"�/�J;�fer��Ѽ[Ƞro���@��gJJ����
�/����y��~��%�i �Y��'����{QrFe��չ8�@C��P o.��5����d�7�nki�!\��m��@C�I���NN����.hp�Gs(��ݠ]����QxW�ؔ�d�;�!���x�;B�~�zУR�Ȗ�j�p�]>�*���c���9��Y)̀"�P[xkAA��J�\���� �l�f^hk���.�Mh�(�s��q�rCe�ƃ��ORo�h.���u��
�~�۲�H�.�t7��lxn'TИ�����2.����[��X���xSB���lG&��7����Љ�y��p�n�ꂿsv����
Ӯ�Gi���V���^:F.R1\O��ɫ�]��{٫,E:NN�Ǖ�Q���Oʥ�f�����ǅ�Ҡ洽39c�zeG�$�B�F�:��	��u��|���%e8�����(�с8Q-�����2��7�X�| ����e_�f�-�U�hHe����`6����]ގ�$j_,�����4���fТ�y|�1�,����R~��l�C����Ba�}��&"�W ����_��)r~��u�t@o�c��3��rJ`���`��^����a�<:��Ȕ�Kq*�2�tɹR �6>�oD��:�frս�:�=�-c�m�(�=�{R�N	K�JD��5�S���g������w:_�"'4Z�_�׌�I��z~�$��;�]H����Qx���)~�T[���Q��<��Q���acգf���JT}�~�.��\�y-ؗ�(��':�L�v�
�o{���(���K�j%�M�+�]��%ީ9� C/r�5V~C� I6X�D�tT�&K�pE*�YI����ُ�K�a��?��7q�T��k�P{Y��V�5�"
є2`�t;��O`��p�
N{�\	�*a����+k��{ �Y��x���z�	o�虊+��G-O��\��������P~<Z*ZE3%:.6a�����K�gM2�|�`�IV0&�%��g�#�ݐ���$�1�������0�CdE�+[E1�{�h�O��{˗��e���q8R ���G$^�Յ��J�`�ꆿ���U#��z��.�^w�R�A����N ��;AE��~2{B,�h�+Dj��B�������Q!CO�q<#�>����F�JG�I��������'�HE����,/&�K�9g(j[�7�6�2�/f=�������b+��#e|�ʃE������,�_"؛S�2�#%U)���7�k�ke��_G��ڇCÌI`ia�j���4v���QO�?Z�OJ�vq*��&�K��K/Lx�J�ћ�������N�h=�+dD_����`�Q@&�Ŏ@T�b82��Gwu�PM��u��W̅U�6�&<���iK��7?H�����J�u��^k�����1K�;��^HNȜ�i�$�3U��J�F��)���C����Dc4J���ڻ^qمO�ࠊXף/>S`�z�Hw�d��Fp���wv7�ն�%�	��R�>�gMyu����1Y�H�I��]?!H����ttgV��mV��)�����w�� ��4���Y�ǧ��4Q�����Ӕm��-G�Kw(��"w�p����D�	�WJ=xR%3��AzKa�X��V�����`j�d��By$��H{���5Rr#i���&0�pK�K�Y�H�G�a6���{��{�.�3����׹��2����nrkF@�U��3%H:D��^�Y9����ᏛuR2:)V�W?pJ����iǡ*�-R����Q�cx>*^�R�[��fl�캙v�5*7]e���ȓX`&K�"M%��[*��)�%��V���Fo���0S/��0]�"6� ��(L"��^3V��*-JJ�v)���x����Z$��Ïr)����<��g���w[ъ� ��tx�"y���\-�Wi�V�K!�z��m�1h�����H��-==d�w(�Y��E~��-V@�^�QAً�Cks����X��V
���%j��w�8�;1��,�ș�ɣڛk����uNӂieY��4�qj7l�i8'��Z�"m��h�.14'�v���*E�|�ҭX�b�o����SA���014� �Q)o�͒I��U���ź"��#1tc�D�e�{�I	f���K���n��.��8a/b�Z��*AY����{A/(�ºLK�G�7����7t��e����tι�3 E@Y�a�^��Wn�dI�;�߳��i��x.�lUŦ�N )K�Kw.��I�2I�Q�$�/��~��`CǴI/GQ5��W��:�4i�DZ]��q����e}�;?�_׎�g��r�0���Ờ�QQ��T�:+!@�N�5��l�4<�kf����ZWi[NS� �L���������%
�G`�����B�=I���[0O��?��$����� ��V�����1x�e�Jy}��;%j����yl��y�ݤ�7�3��遙JzFBa�� ���|�]�7*����#�=l9>QodT\#�<�S�<|��h��kCu���Tm!���|3�P��H��~jeh�!>9.�Ӭd���Z�mWM��"�ڗ9�y�$�0Þ�g1�T���rLw���#������2�ϥ�A��̇^8ȵ�{�gT�,q�ɇq#��ݹ�*eW"����ca;h�"kq�g�]b{��K?>2�;��;>ު�(@Z+LWd�/�V�qgcV�m�i�,�/9�85��"�䶎L\�ʄ�&��5ї�죌�c�6J����"C.nv��y��KfocY%;���4�e��$���DV�S͆uĲ�~��c��eլ���1aZ�.�w�:�9-$��h۲0�R�"Lk,7�x����;/D�lZ��t�I8x��O	����F2�{��gRnT�fg�&q���HH	�6\[YŒ�����oa�L�Tm��q�8�-�P��M�R��`�YR�ZH�� ��_jC��{������d�ଶ��S�^�U���A;,\Pg��<�+ՠ]�����F�p0���G=*>;p#��Jz�{�qN|	���X��Z��P�s;V���^����
��@!�s����5�i�e���{�ك0�;`�׼�	<G����j֐dX_'y�Lӵt�n#���}���'�jy��Mj����+���2K��G��`9��	R�N63�ew>&Aj���cpp�%�K(���a}�;-��������/���`�E��st�T.]T��*��v3��;ǀ�ʊ&2r$-����SB�o��j]+?�nE�1]�E,�EgE-��2�$�ܸH���t��~��E���-���*0}A���(n�l6^�S3���rP�Js�yN�M�(�5ͩ�c��Z����<	�LTL̷ǘ?ts�m�߼
���t�g�Zg0��M��u]��Q�i��uY�J�6���ی>�����xz�\�"Ͽ����*S0�x6/�A��]C1ŝvW V�.c{,i��V�����/J�_��q�Wh��8�ǣ��+QF�2�h�����4-f	s��b\�ӠfxY0H��c��b���_����s���Y�|'O�Y��^�k��|d��ے�8��vo'B�7v�S�[�de�A>^�2Q�-ԟ�BE{'g��p���*r]n��L��m��%�K���p095tN+,~�W�yd� �M( �E�kl+P�ӠpƵ��l�2n��j�Sa ��X�j/���*
�6���D�t�4ٍ:��	�f�����w�u����y��-!R�y�o:{�-�*,���h Z�VA�/Ɣ�ْ�݉\�ݕ�Iӧ�L�������]Qv6��P�����4�~�p)�@??�i���
+bm���i���8��i	��7��Jk������@�([9R�U��EÚU�<�Ev�?f��O��5�$���\0kc�P������RH�Q���e��2���3�f
�3�[���d�x�3kzbu�&�`�z�;w�U2p��~��	d6֘8���-�G02��"f����<���[��ۉ�6���pB�1�"茩�J�x��w�i���gh=�y��E��4n�8����"�(��Q���N��>��Mi���I��ŉ?��Q�t�c�����#^���M�q�K��i��9�v��yT"�0�1��0�l���P���}�alf1��,���%�V�{xf�fy��3��:2K[%sQ�l g��m_aو��,q2	��E-a�5w0p�i�皤߈�ʁt���2�P�_��E3Q����=O���w�r\ y�(s���*�-JJld]�Ӹ*��e��Y�#���T�fc[+�;H�i[�"(�A�z;�����=�3����<�S�����W�Qޛ�O��φ�QQ�)m�3����#��i0��3�������e�Y ����x��S��u�}�.������}i�@u�.����ʜ�ɥ�C�������bz�B^�T,d`�e87oX����;���P�`�}�ӗ _�W���
�
d��W�>�Akv䚢(�8�0�YF��k*�,mHCb�� !e)hX8H���l��R�TO���dxL��;�Zżp�N��W�I��
YJ~R0�٘���B�� 
$���Z�&�0���WY1=R'ۃ1�j�9�A�u��;�瑨�d[NƂ��IqL���.j�ӌ�8�5���[���=t���S��%����	&�5�陿Z����*{����reu��M?�`��r�l�KB��7.c��#�T��@�ҵL;���u��mK�sy/�n��&`����R�@�V������+<w���lb�Z�B<�{Di�z��a{o��bЃy�TG��o[��W]�f]��yc5�ϩ:�.h��'O���*��濫�ɗ����|��]��>���u$��zH�Uû+q��t�M�����Z��&,>��+y^��^r��d��N���n9M�
����.Y":"�z��vn}������<�-��b�v���ݸ"ҏ%���d����qvx8���ҬK�/�Nx8�t�\sOMT��ȼ��mͱ`�A�O�I�7�6�,W��MW1~�_��U*��'�zq�`w���nS
	Ӿ#G�'�y?V%��D�@%R�}���|Qz�^	A�9
�uP��z\$�����t����o	$	��5�:�MTx}�:AjZݨ�x��<xss��k4�Nz�o�j��@O��J���_R�l�җVXb	R,�,M�ڌ�WAI\��514V��ԫ��`%ˋ?��z�i@4�*��"�=|(�+4���M�[�$W�����s�A�ЬYY��W�L�3��&׵�K7�1@���K�牲�iA�{_f�ϣx}��9��?YϜ6G�3Db�P+ю�k>��m(i��s܎r}t4����  ��С��ʣ)<�|��6�=���v/|�!�zү��_EKVܠ'0��,v|Oy��9���`�����j5����)�h�ȏ�����BL�NȈ[�m�j����I���d���y�J�g*]Elڧ`�J��w^8�6��qb��DMm���eg�CB������|�z@h}���d��1�K��B\HSUP��J�\�u:/�P��6Ґd���gf���Mȧ/iO4sz��Oa���0���r �r���[l���[��eϋ�*��m$^N1��5�|�7��L0�c曬�r.���6x�\mh��d�`�#���O��
�������r|zo�?\���:�-gPo�0B�.����^�������.kuH�7hzSV���;������Y�����h��;"�{?��)�?%����!��p~�>X�� [`�@�L�8���PY:�V>j�:�̈́N�*���2���i�ގ�KT�,i��(4,�ʡ�H��Mo�k۹d�` �"�(c�c{���Z�.��[�g6-�H=��ΐ�U
w��k�)n#;+�����Y%}`u�9T�'���GMp�C��I�i����֘�^
ޝ�|j��~�F$ӫ�+v5�O�H�\���>*�7Çꇠ�@\H�@F�],[��폯��I�6��+M=�K��� �~)u�{x�]hJ�-!���=b�7[��ܮBaF3V��'��j�6�L�Sa�qj���y�Sk�KMR��,S�ȿ�oe,˙��ur����Q�Q8ǆ>��T
�G��L(��Ơ���h�>ci([F�~$qڢ��#PC���b���S���Ê�M���Ϟ��H��u{�VS�$!0�q�T/�mԭ����A�� :9]Z����K�N��3��Т묘���(��#Co�E�h�Ǻ$��u�H�7-�yy&��d��=fM^�*�R��#ϻ7MJض2 ,��e(�@/mz�Ϋ�iJ{��i�+�n�f�q=_�X@��9t�I���^�M+���������2Ȓ��~5#7g�hENNDy�X�Ey�.��Q|t�j��B�������g��E&Hr��H>u1�#�ن�ܷr����s7������.�.���$s`8M{5fx���0�捼l�Iw�^�r�������Ì�b�=�"�"�2z����S5G���ڧ5�3���TvݝY�.]R�O� �q�x	���~.�o���z�/��M=2��Kb"(�$G��Ú�$U�4L=��J�L�Ia��LÀ��71�h,�i7C ����Q�k8��.�Z�B΄]���ࣂE��:�H��e�� ���7n�:z�%k���p��~�6�+(��3~C\�*>�% Hu� :��3��Ϭ�$��bOf�j�߲�{5����h�N×�o^�X��G/ᑐ�D���>�P2��XR���EЪ�b��C�'�S:�v����vkY�HDUK7�x���a�)Ϊ~�v@ev�G��x�{3����Y�J��������t9�݅KL���_�0��;��n*x���]��(B-�B�� �rī��NO��f�d+P"��(@��#;n�f^�$	�3湂��3�t��=�Q��v�(�D�����;O`)�{�/��D�m�̜=I� ����O@�i٩�ᘫ���6��c���$E������ .,��y�2s?�X��h�n�o�#V)�ѩa��Q��z���湈�K�8ӑ�s��7�IȾb?�����ȍSk�.UTg��(3�.�ܧo����Y��h��F��b�s/�+����=�^�i�w6���~�䍯�OJU����]mB���>�Ĥ<�-�by�k�l��e��#O���mRS���xͷ��J���++� .�hk�%Q�s]c��TF���_΀	jZ2��(y��ၲ��nT!�uQ�ê:�os.���G��6
�b��t)����� C�h���Bޑ8-�� ×O��v���dv�ԏ�q{Q����,�Ҍ5S]�_���IyCr�qT��1�����ֽ����?�Z����~܎2S(��n۪�U��|9����2�XA�!�qAWh �T���(ݧ'��b�C�B)*���=`�?H������=+��F��x������t�!��WdF��a08�Z�BT8���[���&w�)d�s�j?��"v|��	�b�]Z�vF�k3�Uw��s8�#{J�4$���b�0�jk�q)���1釩ct�^'^�+���N��`;43��ġ��h�~YU���Ϭ�+0s�d�oܐQ�����A����|��/?�"Q8�{�]d���G�?c���� �s�H]��L� I7ż-����Of"�<�\c�\Yj͝Q�"yˬї�+,l��U��48�ˇeYL$�����¦F��S�(�ۃ"�W��E�s׿��H����La~�f[3?vF˻�֔uk�h�~'%]���~�C��N+��[�,y*]v%�Ձ��JH	��!��_������)p�=ߕ:>�ч,;��_\����Q�-a��a4j��D*�Y}�El��Q`9,v �`Ss�/*s��s/��`�(�0I�jz��Zϋ���q�m��3�O}id�E�2�+��]V��a��۶��N��G�1�}�b�,N��~|]kDa���CԁA��7ӌ�U��P����r��,Q�j�_tB�"�B^�M�hNҴ��<5���w�j�}�L�{m�\�0rO�]��d۬ld�����&���S'4<��9��i^�y��.������c��Wv�À]�gkM�!Z!^E_"#U�]�UyE:�K���V��b��0���V�%�A�L�Uf���"�N�4x����V��j%�g���݇���a]��0�nQ��v?!x�#��T����5�<�gV�ʃ���{���䉪�l^�ao�_.�I���X���;�RX= �����gHd����X"�^��5;."p�HЫ�����z6�4J���0�W��>͎dS,7XS���L���f2�vM3�sL\�)*xtħz���'�_�M3Z���!�rbR�T7�-^%�1r���f��-��P��k�ǜ��gFn�,9�q[�5u�̊Y�;y��K��ve���l�u<�2X�����)�4�G��|��t���7$�mHHO%�-'��_�F<��ه_���W�c��fIs�<�V/��9[�)K4:��`*�$�w� ׅM���������\�'��<m\�����.�/�!Ѣ�r��J2촅�N��ze��e�o,'*�B�9.B���$�S���%����D�{?�	{!���^����{w\�>����ʔuW�v����F�F�sm��<�z�D�{���UJ��1�lwJA�A{E�����哔�d~T�H<�@h�jVR�� :���BA��	DYm���P��������~�r���7n!G�R����Kfv�]�m����������m�j�JW?�~#ю# �+ϓA�u_ڍ�[�Ⱦk�̲��G�F��?E���_���(����m�$؎?�ZaZ�y��zN�T�a��to#�3���Ж�%�ξ�.a~�MR�`��b����z�:����+�N�8��(�����P�j��;��C��KH�E68��h�~���J�_��p:�u��h��ho�:��A'�3~#���v��`�KF���z�gv��CMa��3݇�FYv���+5��5��g�8�'��w<������R)��,P�5�8���떚-�l�ďT���F���Ӫt;wj���WS/読\�v�v�>�=}>E'~�7���bԍ��XV8B���#Hλ��V����O�C^��T��;��Aȕ���ޯ�:�P�����"�DR����I稽���e��I~�'"�$����4�D�����"�h�54R��FK��s����E�T�9���d.�N�N���wT�Dπ�(V�Nym'������'�\��l���V��bJ�D�D�w�7G8N0�8����G��e@Gv	Y�"�>�ޣ9�W���6!})qk��� �zp��i؟!����]�#�{A�F������3���gߒ�Q&z�d���:[�y�l� �8j ��>d�P��Bi;n�Y�B��D2x_�`���.�uT�=$}� c�un�B�K���� �$	4uV��3W��ٴe�\{����(�fdk��**�� ��A�d��O��u�S"�F�ʲ��Eɿt��m����"��}+�:!f`Ct=��E*��4GgC�ո��i�2=����=���:�D�kl�=Ts���s se�G]�pJ��d�8��˧gA�r�qb��1+���>В>���WW�,������������������!�ǂIp}Mŗ؋�W�K	��:��^��=�P9���07���N?"h���rb��s$D���H��އ��B����6��B�JE�x��y���J�o���l��&	�\[�^������������
��2I��	��|����o�!��_��Eζ��1���텖?�w�7F7�pi��L�3�]��W\'��[��ָ���x,#R�[hKC��W�J�ɗa)MU[<��Ĕ�S\��&�J7����(�u�����-�OTjv��]�Z��;Q��U��?Ӟ����݌_��
���,��ql��~�X�p��������Ҕ@�������#��T���1.�8c��NW����α(w-��󺆊T��JF�6hR��!������7�_v�9B�8^"����v0nI���K�4���9�ʠ�����AU�t| �A����\
��pњv3im�I�aQj��0=�� G�o7E�+G�NX�#v*j�z�_4�39@Q�v��C��P���p�Zz���@�ZR�o����8ۮݘᐂ�K�[z��t��V�M`	�xX����A6J�x�ò�v��F��<�<pp��f��f
u�e��7�UpP��J���~�݀d�v����,�V�@��2������������:�u�od���+E���*�����m:�s4�s� o�{p�YYv�<ۇ8o>Tl��Ł��p��^�e��Pq�g�c_��9�9��&RսeB/}�-y�Q�¬t��UZ��A���ޤ�R���ʋ�w����eG)�|Zsua����A:��e�˻�G��m��z5kʼR5���
���#Ċ�4�.��񝝅W��׏Et�����F&��ե�0M���@>#$�����}䨭kp�+l0��'e4��y.�0��+	�QpBْ��,O�c,<b��#e4�:�m�`�B�0�_��5�ߺ��<��� T��������MZ�/�BjR��g���-���4���4��N�Z# ]J�H�IihP����+��z��S��xI ;E�O�+�	~h�q��|��^�.*^@�1�Q���y՟-��|M���`����%XW"�[`��T�� g���k���~6�w$������Uۈ������m߳k39V<LQ���B��|cs�v��n�$2H�˂,�����DK<i�*,϶8��K�M�"iN����(�q	_Cƕ��O�T�Ͽҟ��
����o��u=B��n�>9��$p3��Ly/P�][I�3�<a��{�/��}� 8:��Ň˚�C?wV���\��4�ʕ���ں�[�p���݋k�	v~���^7��W��	�!/�M�.̾�����)_7�|�UAUF9@�{�֐��,Â�}&�%b��;�#�k��pE"�H�í\1�3�F�^�B���bl�DDh� �s7�z��Q>�Kg����ZT wڍ�S+�j�,�~�3�lG�>�������cI���ҷ���w	�b��s�=�	��G�E'x4;���bT.�[���d��Hd�i���-|����W��U�@�	<}�	�<�S+�ax�Bi�6�C����tF�ݟ��fy#��0��`����_.d�|�5)Sp���K�2ew��G��/��u�\�m��r��ǭd&���i{�ޮ_��^�"s�����]��	(b�ml�8E�V6���(m/�S��%���t���m٘���/�SN���"�Ot��g����5�b�$�9B����`�Z>���V'����v��tj1u��|޸l�6���NQ� ���J;����C�^��*݌+�V$#��M@�h��߮��E~�`e�ӿ��������e'=���Y��.���8��U�t�tD6|F���c�aw�w2x6ϊ��+��f/;�HͲ��t=C�C��#,����\� ��}A�A��h}/G:�����tx�$�e,��"���pe�1�Q�+
��HN3̰6�(b�ԜS?�Ս�L�c�H�����c�HMx�W	����}\T�� �JU�h������1Ao����a�&{r +��~"g#�����Pk�����I�Mo�/&����Z0����^-�/�G���*��9w`�k� O�Y/@g����_��������U~ j+\č/oNҀ@C�:(��r�0����F������~��gƒ��(8Q��3����8(��ڰ�<@%V�	�G���B����wPh6n��Z�dO��s���6t�V~��U8���l$Q���3@,�9'�AH)��l��'^� �
}��ֺ�u���'��'�k /�����:�%�+b����K���]2@���2>[��~!����P�kh�M�BZ4܈�1(t�O/0���N��f�R<g[侬�x���:��E8R�3iT�� |Mڑx�b�8	%n7�_�x�Ա,=WȨ����U����������R�=�d"J�$7��M��93_�����ޞ�l��KE%/�\�p�X�N�"V�}'�{Fpq�Q������>X�݁�h����vQ������9����3G���@��1h�i,����슖��"#�l�_-o��Jhx�Y�`��g��Q9nD�*Cp��z�����۱M	8�GV�&E�k��{qv���E�y��~���p��Pc �y>B>�`o�.X��$Ն\~3u_/��=��Gy=��;��ʳzC���3�E�_���I�\���
�:=�{���S��G �C�T�љ�v/�1p+�2�9K�K~:r�T�js�|�p4�H���`�&���i�G�$��U��7�}�^�t�̔K�^z�R�#���)�����Cbx��T�l���x^�����ME���:������X�Վmx�ʥ�hD�B��j�"<�̷��xNe���K4������מ0���˻�T�ٺ���,U�?�c�nG	SCI�a\��i�=�lNx�c�m-�5��J����ݼ�ن��C,�H8��Nk[O��j�Q��2�4@B_��v�-�����-)(K���X������(�J*�F�?G>��M�$�ARQy���M�A���
�~���;bg>쾸�ۄCWrh��ʚ�ā���{`��#���$����|-{������1A'8n�n���V�V5��ZG7�:NL���s���5�!�M�#��V��g���Q{�L�S�<�s6X�F\�$/��,���mL�L�]R3J]*ǐS�b�H��@��0�:(�A�>Gc@����;ٮM%ҕ��*��چQ�k���1�qK��>��|l���kw��{Q�����t��X-�!=���j���lm�5�@<Qs�m�5��Z���/�3�Ј��d�3� Z�3֔I�#t���S�]�,��:m���	��"�;O#]��z���	�n��Dœ�YR3J��*�-ݥ�0�T�[P!)@��(j\4�>5��
¦2��v
���K�N�"�=|+21<�i�&��oepz��PPӅѠ�مrFi�4 ���:���ψ���Ƶ0d w	yk�����>E����O�g�&�j��v���F���#
=4�?��X�$�7y�#NaNg�r�Җ�'��]�x�� �'�$���B!�0<��Y���_E�=����Yr&���.Z�\?����@�U:�rLw�%�3�z��@�F�7�&�0���b�,���^�2����G�
���?�$$��.Ͷ�*~��|�p]�[)]�}�e��oZ�{�;G=\I���ä�g�Ɍ�����5A�o,}�pW�l�B"z��y��<B�����Z$YU�����/��,#d�ɥ��������WC�����N�~%wd	l��&�m�o�{x�06�	1ul�@,�b�n�	��4��(n*#�Ze��Ռ]�F�AaSe�=؞����EƘ˒I�W�CeS5�M̃B��h�e-���%_}4��x���sw��C�9���n%y����c�1
��z�b�E�3}4=/|�D[�:�i(f���[:��Ϫ����Z��P�� �Ʈ���-1�(1V�
�}9�t��W��Y��.�"�QL����.�� �B(M>��{`�dfdno�oʻ�2��������yNP��_n�c�"�?Ԣӯ	�<W���b�e��߭���	蓠Þ��h�!�7��W��%4cY���\h�E�u���u�*t�}�M��[5���qI�[mW��tyV��u����CW�*a^�/�c�=�(�IN�8��b�u�Z��7��4â޾�R�?�e�e�{Y���T�Je�v���!� �+R��;?��������6�,n�]m�S|���m��ȥZE��obƞ��Xb����n{� .K �J$Xx�����0��"
Ke��̅�2��1��lx1��W��z���\]ƤD�d�s:��«\g#�-�<�Ү'���'g��Cg%�ol�*�c�c��7T��7W�$� �l�����?�$����X����᳋�Х` )�Īv�ڳ�xExۃ��f*�E�~x�
�+����\q�H��{�P�_W<�=�[f��a� o�["Ҁ!�7��e� ����(3<#��Jze��Pn�h���D�_��e�Pj=������3��#JR��g�4�l��P�gZ=�;��J��eԨ��������>	�P�m���"�o�+9�#��mF�oH�KڵS-�eI��t��V�tj{A���*���G��uϢ64g�t&�K\�k�Q[�N��������Q�=�,J�\�e�	?�b:�o�÷�Kw�RZ��ZR	����5�t2����%��Kx�M.MT������La�hF�\�e0^�k���z��Zn�I��5��s��lXH�Fag$0꺟nAQ��)��t����e}G*ai^��}T��Lm��'��J�*�o[{b��O�}�(���!����[�h� j��M
!h2�K$�;;T|��x�� �jd�>��yH �иw36rJ�G8ਸ਼z�M6E�"RDxHDt[tb+���cauO��3a�W���?�{�*��AJ��XH������ Vj���#0t�)�s�8k�u�s����u�4�9[j��~Ę�o�vՇ�"���J�A]����/��FP"�+�T(���*Վ(h�E�3�܆�6�x��Z�]1]���٦]ݪ~.J7q|7^j�S��a�2�~����\�D���&G����,�[���RB��R��oa�R��쑢������,%�ᒻ/1R�v��?�����I�i�򗳭'����{0=�y�5�Fi�5�6=W~����o0!�ԏ���։�h4 �zN,o�I#̰����Tig�8�s��CI1aPʳ|�pW�X�/걪p�>�#�0��x"}�S��$_|���]M�z�0+L��C�
���3�J���n������'άV<�2a-�G5`o:T˖e�y��T��NCp_�<��V !h�����?N�y:��
1�f]+�s����ۊS��,nL�n��vF�z=3h���8�!Vs�� -�ҵ����P2��q�U���u��>�<�4�ϒ!+��&�����a^���Pl��b䚬����_��ȣ������X�^쑬+-)s�05���q��{�]�ŧ<i_�>LZB[��_���u�C�x��C�M~�Y`�
��h���o5��)��A^���8�*A�i-k:㬦�N�֧�ޏ�"�jm|S��6hB�~X"�~��蹛��Te��w�>�P@�L�/Vu(3B�YP� T��I(�z0�7IP�{��3�?�3}`gt4�X���B��t%���)C����Z�m�t*8Ҧx@
�R&�Κ�P&X��/�w�(�g�VK�����e�>eJ�Z[���}?�'F�<�(:�u��m����m �W��W��ū��;Og����K\���c�x^MCDrp���*��̅��FjMe6�4[�Bfn����َ���&��nZa^��x�Y99�l�?����o7�:�jY�&nB�����WBx냂-w���8�T����I5���cNR����^ze�I�߄o��.�>O�z�s�Nbqp��rJ6�e���ͫ���^H�̹�>��$?�b���Q���D5NK�W֢��W��"�����X�����2������hM(Nay2;/]�ڱ�����,ށĎ�X��Ē����
��M�k��6�����~��K<LV�]^S�*19���G�����k�<T�]��VsuMuO�h��n����	��cF�vz�<Rƿ5��EPGג6(Y�Jl$�mVG�s�o����ʡҐ�}f� i�G�b�)t,�.~N8���4�|)C��a	݀v�z���`�DD����e��4b.���������o�Je���ǋe8�o�#��,U�rz~z������ؚ�8!bѠ>�AU�X�	��y�a�Q�"�L���Bo��C�ICp��=b�;O�$$H<�Ŧk�z�d�\+���}M�M�]�p�c59����娅�	X���t*�=��MbA�֎�o���|2$��XRM�A�<v��L(h�Z(lx�w&�>��o�3V�x&Y_�E�B��K�Ac���I���v�!$����P u4�V��KXy�̈́�Hix~�!W����UAN�����pR��򛨇���?���ڣ�O��Xԟ��+�km�:!sޥ�n<.��4q�%��eo��HM���������§ P2m8��^z/�j�v��R�U�ڟr��F���!z�5���-= ������i1��@�1�Iƃ��b��x���m�N�G��L��lhA@� p}i�U�� ���[<�$�r@m��Ժ�K���>�c�)�U:#��e=�}{Z4�T&�BD=W����<���'�&���/W�Ea`���@��B���5�>��Uv ��22ߡ��G膊_s����kd���Wa�u�ލDD��̒d7n��9�bxr�5$R��{�b�/��]�c�gh�$M��0gý�3"���Y}����׺КXLZ�T�����2��vU��6����6	^��Z�g���g	�A�Ǖ�_L��k"$��@���]{��V@�^����CNu�nC����3�)�7e��[�zcF�;NMPתa��D�j�<��T\j�ˌ�`�[M�+1�x�K��]~n�z;�l7IZV]r�*�� �O~>̹�?+c�-!l��6Aǋ�{����l	�q���J���9g�xvEi�kł�X��2E&�WԴ�הVM��=S)C&��q����;4��0R���@~k��hߔ�|����8��F�%I��#�i^O��O�vy�,�����z4�|�f�m��冮m����@}�!��/��m !�ŝ -XEzw�H+'E��_�4����R�ե���"�2�Q`Τ?ջ�v��ԁg3�zXj��	 ��ʍ3���x8pZ�t��1���Y{,��w�����Y*���ǵ	��ȶhv�_E6e��[��p���N%aUJUf�Y��,[�:#���\�Y5v���~�:�ob��S�����!�\k���+�V*w�d�K��P����o���$*�����/r��%�=�x!��6����>��~f)~yR@i���zc4��g�e����9rQ�jGJ*��n$�e�liio���
H�b9��9�@�l�#O=��®w���8��'�7����Z0����{�:R�8ꬑ��)n�W�v�笸��$աC =���X9ȕ�TF�+F��-��߂ً�NA�ўo��>|�[��wz�ࡕ�D4���~�-(�����5DY�&�pnZ'#���q���8��Q��UO,�+V�?T����chs����&?ݧ�:X�W0��C�GoEl�
�]�������5\�3� �2��A�So	9�1M��^�P��]�89\����B���j��������bwz�7[k=��Q i�~4�ʑ.�Rf!N���"/hk(�,�I޹�f�Բ�<�N�1�hW���c M��x�`��ͥAJYY��E�bLeq)��6���j �-��:X�ׄ��5p�cH��r�������z
i.g;E��H�HN(k/���P�����ʄ�q-�ĵM��٧C?�Z�u'\��a���o�0��?7��p!
�_��1�`����3��3Gm �K��#�<٠�K�~1ڗ�h��*ř��Xh�XJ��3p�]����a�;k�k}��D7|���,���3���4t�xC�ןw��E�0+@9U�"�~3:r	Q�4"�鮘�.����ື�I_��2��9kע�.�ɦ�=���!���9I���yXN��A��[?I����6m&ll�z>o��]���JU6*��S��A��Q7�t=D"0���LU�T���kK/���8����G��)���I��Q�Ϟ�O�o\�';"�D�Ku��5��m�LE�X�sOz#}��Z�I�p�9)�_�W=J�H���k������凴4�wl�����(���ic��WR�{O=n�Xh��b�ٱ�#�$�(�5_�za��59��BqԽ���޵�i��>,��i����j�	Lc`��~�f������;=�\H:��A�� ��]+y���f��+�ꥈ�L��q0Ɂ$/A�[De�Wf<pc�(��
��d���;'��� ��\��U.߈��q��M#ԣ����r��#|O#���y���K�X���=�H9���}T�f�5ō�06��>��	}��[���P\	�4a:�u�&J�,�Q�x����j\�0٘2�9+`�",-e����#Vtp8�#��'�%.�����fܻr�ڣ��$�� ��z%���U���E��0��V��,-D�"�<O�qd��oe�2��1K�3Ay&���5��{�<��V���o
����摨��96�6e,G��E(�\
��[��]�<^��E�۞SH*�R��N��� �X�Z��Ff	.5�$���}2�IpY;Jh�ݿc^o��p��cgfռXTb{�r	���),w�ߚ��ޠ��뢊l�'%1a�_�8�Qָ�z�L c�.��7�R��nJBTSC0Gf�J��876�[�����9!l�#�`�~�>�����j�{�f�n��,a��u�`��PydW�����)6���ι�K��I��D��©�mW[M��� b������RB���o%���`����Rc��/:�Al�3�J(����=."`Tu*~a�-��X[�Apy���#Z��K��z�݉i�<ob�B�&����Gq)$�f^"*�ڂ;���C�6���3���a���`[;n��C<�DW-
Y1\��R��p�
�
V���#eH�'���4^�_��P^{���h[qӝ�)9˴�>i(��}f?�K�.04�����d�EJ:�Q���N�Y{��/S}� $ii^�FN=��toY|�镓T��7=F˗�4h
R �L��?���U����|^.<�����,�W�6�:�I��;6�����p�u�C Y^��>UV�;��c�j ���O#�LV��9��|�{�U�mk6P�}����kڗ�K!����Y��\�"�DF��ǖfӃo�U��dT��l�,����ә��H��gN�����3�ϣ����	Rh��y���� 3�
���J!JWI�H2�����:J-cר3b,OI����DH'�$�q�7=kx����c�ɴ.8�X'ɭB��_u�?��2�r�>�&%n�6�An�
ӕtqnai̎�V4�l=-�#��'q��w1����%&:^����>���G'O��g��	��tB�"�9.��V������4,:ֽ		�m<pd���%�_���!i@�R�X!M��9�@�5��;<i��+H�ٛw����΍.xz�)~}��p��|�S�D���y�q�b��-u��
���/�;}:S;��������*ꑴ��-i}�92ϹӔ�,L����!.�����#�q��ɚ�-2��~ui�
d%$G�y}�S6�ɶ������x0Ӭ�{X8DEx ӗ�f�.E\���n)a�m;���?~ܷ*�%[M�G����$'q&d�9�T�V4s�8rN��W��|[��QR��I�`k�j�o��YeӉ��=�'_4�� zdYѠEMsf��n��A1�ƍ�����5{^�;��jSNs9��!�àl��	EZ'Y���#s�J��T��Y.�e��ʊKp��ꗘk����Ka\��f��y1.�}���t�2��Vf_��*������3U��ٜ��ۚz`�Ж�#�ޔQ�Gb腵C�l�B���ŭ�<
n�H�"^�`K�/4X�;���q�RS�����W�ӣ�ە���kf���c�,���}DvźC�,�T���	!:�?�H����ͬ��~�����z!�/턉�_H����p��>���k�._�H}�V�JS�yC�QWK �N��4�FY�
8v2�ct�Ӓ褖+��,���p�m�^d�_ڸQ��W3C(ŝ/�Y�kt����b�C&��Ǌ�	펹�JO��补���\\O���4� 75W����9�`o�\	ܾ�J�ޫ��q఻��=��糣Ϣa���8����~�6-6[Uac.wm��efx$����UgL�s���`��\�{<G���&톀�"N��2�~��' 9����X�C§�	R4���!E?E�f6?�E��ݥ9gTH���v�m��;-�ХB�D���_>��)�����%G��bQPO�03���[n���P�M	�i<9�{*'���'>�
�t~q��v�A��ѮAP���l�1m�^�Z���d*�u{�@�|%���}����~��;{���V�1�#7	�ן�H�'
E���u4`�9���)�h����Su�T��t�
m
�QN&�@�p�@\A>"�q�-��n2��b�-ы���Q��#��-�5�Ng��8�Zg�o�c��?��q�ܻR���\�O�ҍxa�� 1ٵ<qlr��G�f���U�K�I.�
br��Z�����E�:��_��i%��xf����q�����}��Mx�2
�������)�i������ ���E��6���\~Ӹ��	p���Su˧�}~Ei�����`�����t�t�k�����
�듹��wI��!!l6r5ű@ǌ|L:N�M��KߦD��F�(Q|ai�����	>b���`���x�_�%��	��m���>�LEH�i��*�Up`�(�����ǫɜگ�/`�H��
}͉�q�hQqd�M�)��	H:Nq�����[�Iy�ƶ�Q��T���]|���� v��^h����˺�<,���ԗ.�D��� ���y���+������Bvu��?,i~���pr�)��U�P����T��'�ƥ�,����������+��ϡE(�Z�LCP������' �p�L�}CҀ�bژNB�@h�_�ͯJ��=W)�}Xs��S~"c�Mz#� ���T0�;��H�����S���V�p!���� MF!�����+�#fHwUa6Vb��`�@��f�bx���*���h+z�XJ����(UK�~���]0,l�r�0��T�oRѴ�����7��"�r3Vؓ��W�R�zŁ�Vm;o��_ᛩ�z�Uat�o�%"�1��<ݤ�19`��(�_܉AB�Ը���|�M��p�5�*��IMG:�B��ZD�x�ɫ^���Q�9�f;���A��k�Nr��9�Ux���w��=w\�k��U��'{Z�#)yU�5[��c�k['	��,�ͿY�E��k&s�Xj9'rL�~��E��h�dO���w!�����lv�m��}ܪ�d-�$E�7�kAC��J��3팾�.�H)��vé�
ZX�3EE��V��~��1�`c��fX'"��i
����E5��������ԅ#�}�g����0���Kl�6Ӹ<e_�	�t�:x� �����'���#�n��Ɉ �6�ܼ��GZt���P/��P�c���܋�@R����(�+9[H�lQ��% ��c@#~.$����az��{�<ȶ^�Λ��z�ӥ|�G�� ia�9/���b��`<�cP+��G/5��n���$�i�S�1X�ϸ��A4]Z���JR�%h����0��K��9�G���<�n������[����N��2�(���_O�=�S6oۘC�]_H~%蓑��t������N ��[�B�Ǣ���4_�}�~��VDT_��~��ؔ�V���
X�?B@Ӟ{\�l�J=J.��Ԃ�
jp����t�;<�,�!iH�)�X���AAab��w�}9aL��[�Z&㢳���μ�>�1��X��ѿ���J�ݰ����W��V��.~��I,I[druW�&�N�AE�����j�B�;���itm���֩lLEU��׽z���YV9ʔf�+5�9կ�3��}.?c�A0�v�� B�{���Fx-��\�nTU�Ы�tD���`񕓁pbk���!��w�0�퉤�;9�Ћ��)���6�w��t{���Er�O�\�-����(rcj���6U��Tcg#��Ԫd��1�����I�R#n�%�=8Pi��H �o/��M'j4�DI��s�Oc�MN�.s�|��>g�}�o�v�F�F��)�+�.j*}��R�M�d�A��R���{N�6w�m��KM��6����_����z ���Smt��v'Ufr�o��г������W��<TI�=��򬄫�>�wd�U�5���-�d̕i��*32Qgϼw�Z����fS��1�RM�a-�Z�3�o�ak�o>��Q����Tj�����ڴ(�g-ڮϽ�3Gn���ۆYo$	i%i_ߧ���ְP�1՟j�T��u�����1�>��V8�[I�|���O��v�)
����Э�zuB���5��D�t \>av�=��8��B�:�ݞ̕�_.��E�����uv>Ӻ#+/Z#RR�o�-2b3찣�;Lnۀ�e���=�U����n<�c��=e-z�����ϸh�d��o���,$�A�Ō.ѠC���Y^�l�D-2׷�Q5	컇R�n��$@?� J�\Z8i6��ĺA�4��zG��x+V�����II���h���z0~��f���d�ˆ��h��1�)��z���v�m�	NEn������q�_X��	6&a���5 �^m�Q�RjhX�処],)�4�\a&)�3�APF�*�V���[ ��g��8*0Q�s��%ǵ+B4eղH��Ɵ׬mYI��q�^K�i-�j}����U
9����]͋'bg�<����Ry8��턭Y1܇��G���HN><��l�V�pnf�Bi�ju|܁��?�����~!9x6-ʘ�z��Śx�\�f��e�����47��E�Vs
�����:����#� ���d�j�"CD
�Co�1�+��ho���N&��T�jx��[���35���|C�vE}��9�T*J�Rlpҗ>�X���~=��6V��˳A�am͝����5 �\:Ы{���\W��&a����`�SP�ǹ_O��f���įb��m7�8~���K�Lq�j��^F�F-�CQ�)�����i���������=,+#���E-cSg���)���I��[h���uc�5	Z���Y�ڪ�`��H�]��85�M`��v��"C��[�`W��hE��D'�a�FF#2��^�mS�oO��a�=ݛ�
��7�|\n�꣠� �h��������R������If��������5�(�����}Yi��ԐܠN��)��m>�NJ��ӷ6N�����i�+]e[ڶ�ߚt)��\�xb]"$�!f�ݴ��'����,&��,���0�� ��A�٤�*%Upt�A�X��l��β�gN!ŔiE)Ɉrtr��5�!��R	�b�L�~'���v}�3��0��A��������6C����Q��^Q�躰����>3�&J�/�i`�#��h�D0�6��ء=$?�G��:�s�1�r���gR��J��&�+j`d�Z=�J����Л[���e� �f�0�W����]-(���v�]�(&�����"��0��b��ɞ�>���43i�VX��<��=O��Rd5!
$�w@U��5�"^lwBwo;H���@�4�z�]c���s�Ow *�9�z�!�Yl��.��c}�����8�����<����5�`�Ӂ7���1�^��-���E�>��Rms�F��Yr>?;��9W{yц<�� �@� ������eD�[uZr����;����K�=2HӖ�m��z�8���k)�����]�sQ�2 p���B)Z��clD���%��l�t>Jn�_IdZ�@�4M�y6v���h�� ���>����oG5i5T%�f�|^́�al�IƓ����_��.�� Z1A슪ܭ�k�/xS���{��11ҋ���
2A8�v���2��(V�����~!���k�NY�l���do����D���Zج^LIqKhkYJ��
���[�%�8�ފ�X�0!c�.�Tw�^�bR��4�\;i���W&��B�NA{&��h5)��-hVӺd�
���@L������b�l��Ɣ�����"G�%�d!��_ZY�cz����0������n�:6"&|2��!����>���v���)�R-@�?��O�%JD���r�uf?P�Vׄ\�t�]�qa{�f���kw�����Ȋ�y�j$��.T�? k�%���l��+��[�,�?��Î �k�f�x��TD����K��L �Ӆ;=�ywɸ^�Z���aM9>��գp��[�Y�h|M#q�'���8}��/m�Vb��n5���nڂ��bY��������+�n���I=�}<�����r6K/��[�$�U��9��D<�D�Ǌ�|X}�ϒ�8�vT��@�hW�TF�?�� ����a4q�I�>�Y�����P{���eAB���'�&�bTp�]]��g�i��m���ݚf�Wo��(��� ��*��T���We����B�V�j�VL����7�"��?�[mb�P�����������ߍ�� �UH!��t�g*k]Rh=��>��TE��ۤ����9dD��@,��qgq����P����yv�BTFv��������ڋR?!&�a=<�W��;�'F�KW�g�q�3�����=G��"��S-ŵ�wG��DF/.G�7w���h��v"�Oa%^�=�[}w���%�v 6���vd,mKK����6i�4ꍕ���?�;���������u{�:�{%���<K���.f5�c���E'�a��o(g6���Umqj{LE:�q�g��j>^W����芕�W!_��ta���U�e���֡� �nl@�q;�v�pH0����\��h���7��OC�M��{R��!Y��2,���IS�k����[~j���yd%YGl�P�{�m��#IY�X[��a����'8*��^��J�ɲ�LWTw��y%յ����y�������i�Wb�lZ;�ݪ>z\bC$�cC	O^jT(@�.����^'8�)��T���� 6�"��2�1��>��O߁K�2l|g�F�_��T�x��`y����9�8N�3��Sxp�#Hv��hQ$���^v�����GO���γ��|��mY��,#=��/�X~Ш@�	g��!��YT"�2dd,�=&2������eF��/O��A�d���b��K�y�u��Ȅ�k/��-8�Tu���] ]01�8�{�����%7fO�.�C��f�n��Ke��j?�E��)׾h���N���7�A����l�.�{ջ��ݶ��6o�f�]�� pj̹���/�|�z~�w�1z.�	�B�Y���rsS,�JpC�śH���`)����N�{�g�oL�Mj�����k�� �f���2d�v�"i�6��O�s@�Z�P�)�m�*Vjїjag����Z`���N�@/1P!�A��� ����-$��H�}�UU�ozSm��q|pNJ:�� ���@�ӳ�c�x��y�G�b̧���H�Un�ϣ�
;@>^�H��&QmO�=/
ߍamh��V��r��VT
�RJ�ϳ�����xi|B�z˨�����N9"3K �.5�	�vPd2��]�L>�vh�9l�����E�v�t� ;�ľh��.�1	� �L����c���#|:��xc�=[Q�a�@��h�c�װ�3�%k@���)�ڝ.���{YT���$0o$Rz���N����X0��;!��֚��FC�t�ms�QM�M�8��m�&��T����ɂ���(�g��8�&l�����zB�	R^ȣ��Ap�s6w'_�6o\�VC9Z���?e�皥�\�	J�l7��{��3���vo]=��7`��1X�p���s��i��Ɋ�2n��ɒO�s+��|��d`n"���O�]��)�l�ׇq=�b�Cױ1Pۿ#kp�Oi]�bC���<���(�zBhb	�����?����m�Bņ@�<R�ئh�>zxd_�j�W�h{vp��:�oy��?,���\��)h%�}�Rt��$k��۴��}cD쳉��6�>�����$�j�4���؈��!��P? �����H�W��c;{7�c�����b����|$�I���f3\�8s�!'H$=��s����������8ܒ����M����%�
��,�	'�_��wx�4���ׂ2�2#�-��2w�{�H���}�|]������a�\�iKm_{���N�Ai�����d��N�5�yiCIN��h]pGr�(��RD�[D_�Y0�ֵo-�����ƏF=�c4G�ձ��a���p�
�;|�qxZi*n�c�(�Yv��W�qɚ�x"��B1������7yxZv-�ү`��
p>"�iEw��1y�s���h����<D�b���S��ou;Ͳ'.��F١
�
�b�s��CIQ��GV��^8<fM�����ڪv^��@H~Y�[b䨵Fk�k �� j��}ܯD��8���o#��� ӹ~�V�
눀l�)�L�MU�V1���5K=���h$�8%��Jȉm��1�&�0uV{�b�G��?�����E�Α7�Pw�,	�<|�M�.Z'�<
aK������v.��'b��c��Ѱ��~�r}�D�����7b!߳�)d�ZtW�=ߟ�DÓ	CK�߿�����tO����0<��̀���w���{E�3��ޒ"����0����J0��]��vt�Z=d��ʹ������@1S���B��<p�-�G�o�+��s�+1ʵ�O�~Y�ѣzv������Q^}�X�TN�UZ[
�W�]_x�4-Z5i�`:�XwNU�\�^�$1�)����У�Sg0�z[:�p@���a�̄L��lJ&k�Y$�V@EfR�g��SY[�|F����g<G�X4�X�c���ܼf��L��3��N�vns��X�Y^;�B���Ŕ3g>]���\�ț�d�wM���qs7��&�ȼAl`���{^�����u���k��,������8'\�1i�G]�i�+3fF����0�]9�vYЕ���]���_]sP�j����ܲ��J�*������p��������}���y)`B|U�?V�4)�	�E¯IP�GE�%�/楺&sƜT������֘�l�~����/�����J�Q�[4Z��VR�O�PZO~L�5� �R�_�ČS6�ٕYp�L��L���	���O������r���&	���o��Kf�=�������g0���ĥ�;�(Ȉ��by�N�_�\�]�"�΅M�z�� �n�-������P��� _iS�6I�Ƹ�R��9&���%P �
;�U�c�8Y��E����a���Y�	i"3�w���4�T�_��q��p�Y��ȧ_����0�3x��ը�>�p �� �0]�W���!�	���	��Mκ�44��@1��k���7H���Qd�9��a>�[$PĖZt7O���_�"�JV��%�[z�,�b��`�#G��)��i���3X�	���9����.��V���)<�2��a7S{�pzi/#�'[�z��X�)L4�+�SVV�'u�x��l[��9B��ic���a�<��2� 7I��)�ݐ�u3r�j��6B����>�"�_���xTr�t�����)n{e֧�c��s���m�1��(%ه�%�FD���O܃�"3혗�)A��6r�F�v�mv奆=��c���{��Q���p���� ��O���&�ỏ� ��S X��+�����)Y�a��'��j��X����1�#�Q`a�|�"�׈�~��g	��#����M,:Ujl��j����||�I���-�"3���!;���K?�7���^a<5[����%������~�Í�0�^�D���Z4�����ܥ�X�p���L���ōA1����T>90ͺz�_��.���ѫ�8vt=Td�g�t���Hl�-�iq���8��&)~�Rϖ�Ir�l�wZ߱w��X���)-�q�,^j��"�w���PRg��F�Ǣ:��O�����Q8a�S/�)Zg�Y��PK�:�r�ei	��9��8ٓ��O�xb�	��_$��j�=��G&^Ě���,΋�4����RY�L^��T��\��7~��?��J��6o�a���Y�Z�_c�l�@H�?y���7�R�M�����K�m�h����*��m���]���=X1�����@��R�nU � �N�M����Hjy�w�d���^�j�K��^QY=A��� uDKM~�QT�]Ǽ�J�oJ93����]�V�"o��'��?���z�23�x-�Y��/���p�K�{�hvc�>�����#�r����Fr'�c���bN|�P�����"����}���8\Ҏ��w�J�uV����-�Ƅ�{3Z�)%ax�/��ߏ?��Ϡ���
*����.$̤Ue����z�����I�,�",*K���S,j�)=�en�(�2*��J��L@Bh��� s��P7�ʰ�A�{��}�ʰ׌�'(C��`z�tl8������o�ߨ�]�v��ю�`�<cQ?v�5�ʚ�]���fE3k��r�l���洷�`xIf�JzM�Y�W�l�@��.Rse���:+ܨ��^�8Bp��z�K0�^��~d�x�C�"��Vz�
����ъ���v�gV�!7g��?R��l���.�����kT4��TS�-C\%�<��G�	}�~>zz�s FT@���X)B�Ju��|�����M	R(Lj�Fy+ܜ$�vJ	^&��"������FEA�� �lI���D R@>��P
n��&�;��M��=�$�M����
7DˡŤp�"P�\Ap� C�M�5u#�9��6f
5l�%��g5,��_ZP�b�\���'���l� �S��W]SO��?̺��/�p��~��z�
fu|��o%� �����?�F)ż�ޮ�0jbޏ��2BG־N�]�����hV��� �tnV��C-t�Y�8a�j�(nI$W��r1f��B�hX8�duX.��>�nҹ7r`1��Ļ��!%�(��	_FV;e�ŦLءE����|�jy��%�(��>y�������IW����x�i/<P-'�;��c?�2���C�-Kӎ�q�9Q�����zK�9C���z�҂3Wd���1$rw���%��O0�AY�3�J�md9U���8aKD,��(��f}*��؇�A�\�N��+�50C�Q��FW��sK�?1�?���e\I��\|�7�ο�Q&�E��^(x�&��)���.����H'Itc�\���c&�>��0��������m�T�ǁ}�gKFr�B�N��%���0tP�M�*K��(� `U����H#� �>B?�@� b�K��o�"�x6�.������
�o���lNz ��o�E��#����
W	����7�\Ub/Cf�:"c�O�SO�$9�.��d���u���y�-�[�뷩��j疭
~X�D8���_#?@d�ۃ��	��%�p�w�o{�	L��+�9��`{��7_Z��I��*�V�׹�V�(vd��g
<mU[苠�W�� �ܒBhK����ܞ;���+���浄��ۘ�/o�̠lg#^o��XV�9$�D=�t�Q)f���.4�K�/�'���	n\��M��L
|�D~�O�h���Q�a�:A�y
�o�|[�����ٟ�r鑇 Қ?��s�73z$��σvD�*�����3�g�-c�6��@�v�X�E���Ϭ�Zϸ�gO%q+\�6s��/����h�	A��r�>gc`��`�S�?���гjt�9I4O�����~t�w�Q&�i��3�>�<7��&��8���`�S���Ƽp;K�{ٗ��@���cQ�6	�6g/\����K�I"�XݷnG��i�^���׾I�R7C����n/���1*F`(A�5T%��0УW���g>�q�Cq���SF�<P�,��W�V�8���]ȩ�~����Ή"Rp�ɀַ�2f0����8�!w������/�;�-B����P鏏���o��d^�t[.);��%�����[�����J[/N�$I��K�Mn��5����v�@��uK�����2��B����'i*���/D��5���b��������}�A�Î~Tk䭏�<����I�b��` )�!5���Чm��Yz�����;̿��A��^�ywv*�Z��ߕj�`��
���?tvb�������h�D~�D�W4h�A�WO���Bi	s��r�a�~Fg�����|�̔�����D\7.g|�!��Ӹ��T����d�QgbF��xx��w�����z��*��JX��<���f��f�>ґp�ȋe�����%n�g'���7qo´��D;�űF�&&ۆ�Y��1f���4��&�VL�7��Ư�p���V���n��p��#�t@h�(��J���l�%���#�=�2v����[��8W0@�nX��%���2�ơ��~�s��r�豽J�j�����<� ���DJ�+7LsS�^<��ʥ��>rt�E{\���,'�Al�T� �4�lt��KC��Å�AWB&�쀀���s3�-5��k�L5�2�}j���D��I�w�S�y;e6e��Ӎ�e]ɨE�1�u_�,5��L�����������[Ry+;k8r�e�2S��sQ/���T��h#�D�@� ��v�d�;�����b����p�\b	�?r�[���ĎL*5�D��Dr�a�v�W/,eC�� &��{^�;�q'�5ֺ�PF�K�*%��)D���g`�qzM�4љ;�s�1��&��(Ma�ҟ��d�����9���q`�#{R��*y�O��_�/8����;�u����u�NB�f�$�>ŉc�Y�%�ֱ��%�S}��$��=�K��y����%"
*������A�w;�G`-!�Ӯn���6I���ew�w#�i-���%��Rxe�C�1v>V���XȺ9M`>���6 �f,W(#�j���
�ں(7)��M��È(�=�Ɓ���e�Z7�:xﵠLҧ���o���k�X��o�=�f����ں���ɣx��G�\0Yu�嵧-&�/����2��]4s1�'PQ�T�f΅�����0;m��z��#��3j�+��Z�]�ׅ�(u���yR �W�1�I{�h���"�~<�a~PusA�C����F�p��V�����[8�Lij{�_����{�7�L/�Xb�ѷ))���Hױ�Ԭz�����{�M�
]�h��.H���3�����U�)�@������*�=!�0&�"�|h-�P�ﾝ7�!0� ��R���)�\���̵1F��\���V�Iz�F���˶̨)����3�=&g˽`�R������磊��+��aD���P5�$��&���:P�NaO��O��5̽ȉŲӱ�l6�!/uG~�\>$���� �~�aQ�A�ɥ7N�r��vd$P�>Wy����w��=˻�[S��)�Wdз�;���RmsW�"A�tH���E���/�V�9�7�j"\�9,�"? Iͧ�����YF�f!�����#pRU3��Ht�3� #�k��S�IF���E�p�c��Ԧ�Ʋ��%�+b;V��W�u:X�!��Ҝ8�^����t�]�RX�<�~��ul�{�����rLG�]g�� �të(���I����t�D�,��ϻǙ(���rc'�JL���LY���v�����
�b�t�P0(w���^�F��"
~ՋQ�@<��� ���_2`��v�-2m�	���Y)x��W^E�xuH"1"�^j�e�ˍ�'��R���E~=�Ⴠ�#^�$ï4�#�$�|�-@��
�meѽ�;�4�=��+H�O�@B�!>A��(Z$t&İ�����[�Λ��`"���Q���t�ʧ�zږ��
�����l�$|�_%Cx������0р�m4r��B��%ha�D�N>p�����>�?��I���8U"=)9���!`���7 X� �6��� It��A��9�����י���1�4uM�7�z���8��'�/�jTo�y�
��:�c?�x�L �S� ��]��̕:�d��X�"�Tr�<MY�nk��'XJ�K��).`�.�k)�4��+V�����7�#U/I�����E`0�����gL6ԑ��}�%y��5��t���Tz�c1	�pU�����s(ہB� P�x�\w[���l������l\c�l��ʼBOf����po�O����pxd��H�N��Y�dS[BkLr�ۊO�]�Mf7��q�Kxȇ�G�]�����yz�g=I�j����d�3(cy�)&�iN�I ��|e�8�����Y����-p����v��7��$�9���ǹC���JZ��R�2h6���9���"�@zd$�� ��o�ց����MY��	�=��M��bI���^�X�_,!�jn��o䖆Hף��ׅGh��+i�iAT���]�
-,F�8�-P'��КAͽ^��w�
���_�GWO\���B�a��!�����	GT�������=?���N��X<[�쮵��Se��X��,�j��j�Ô��+��`W2�&�,�U]pK���R8��9(��s���<��x�c���d=$p��L��&�E!�X.�'o�eo�8-c�/�9,�.��[�����?��K��!||���*�"���P�
�57�'��L�s��ju�
ِ�D�w�*#]ȅ ��]����&�/����S��m�'*,�o��d��Y3XA�L�'�~w:5&Ї�vJOJb��fR�%*�w#��aJ�eFc4�4�@<�����&�8g[�\qV�d� �u3��G�RV3Ĩ�8 � �
�Ր�F�+��`i���WBK�ދ`��&�]3��J����/�F�{�1�שicJQU�;YH������Ǜ`A�y6,~�b���3��t�^-X� �nd���oa��K�URQ���ς���n�E�)��6���;��˼�w��cXLD_F���.>ڍ�U�5���Qc�v���A��8|�Q�UCR��ߙ	i:��r6�����$Tb-�VV��NzDW~�G����P�i7��A�:ߎ2U��ͩ���{��S#�ڸ�ݨ�l�C�ܷ�80��|2�ȣ���	��U����h�j�>_���:"]���Ki�sH�<�F�&�1p_���
�����-΂N��C���Pr�Y�PܫB$�_L�W�^v8�x��ʒ�'�<�<܀����$����H����9�RʪWA>�r]�;9ᆇeb����˄�CnRƂIH��Kͬ�*���(v�J�jH��#Q��0�_�Ȳ	�Tޔ��0��eƅ�.��$?S֎-z<���ũ̺�R 1i�����l�!K/���,���Դ�������A�������m(s+�|�c��!T�:���}���cX>��5���v��F��2�ԻL����du`B_I]���g����-���L��%DM8��X�V�=���x*���Y���L��#݋�]C�S���H&Һ��y!�gZd������bX;ٛp��g�L��}7�B�G��2P?���jٽ�+<+�G�+��0"/�e����Iפ$�|��ID��V�R.�V�L��ŗ�`�����N���w�ڷ�߀��:<�f����b���\�k0�?�~P�B.�d��kgP>�m�O.d/��G��������6~DsW��w�%Yz��QV�
���3@�R<������)rH�����j8^Qy��׻k�B�ɳ�]d2!Ě_-��]�UwoՑ�+��z�2	t<��z��A<1�m\CPF�F�Y[��z��߇(R߭k�ܢX�[ӝ��uS���֋S2�n:ta>�z~X5!$��Qg��]����4ٺ6f�p�ɘ\�]=�	\Ǯk>������P����:��(V��5;ч��V	n��pQWE�� ��9w\h�('!*����]����+���G%u�MACMx�������\����:dsGC��&ܘZNc�##�j6H���%C��EHSG��x	W�>;v���bS',�i�O��L��d��s$��<S@8� �i���=�.��u���u���1�uCF�>��]������M�.�V)Q�#�Lr���)cvZac=��h}�������H*.�J\Q��6�ώ|��-�Q��zI�	��@���-��9&q�VO.�O��ʓ���J���>F�AC���pNa%��ԩ�ތ�D�Y�1Ƚ�Py�ɥ�Xwwg�q�b��J6KX���8@Z�l[�s��<�bCl4J��Jﵮ�i�(�˾]��{bG)l&���3a�B1�Y�=�6����7�(���ݤ��]B���)[���\�ϽJ����Wt���]+>����PC~�)z�U� t���"4*�8�)���}$ur�1G�8m.�i���r���Ƕ������V�5MօS�VO����J5��{�>�%��0Œ�V�q �ښiG(�3I��͉��K���p�`)��h6��*qϴVt%]�3b:1q�������aG�6����56o�uJ|e�+�˻�9=�o�[wǛ�r)i�v�\����E�V�p�C�z̦{�r�%��2b�e$vcL�r��{�P���[1��qk"d�VF@K�ug$�Ms��qFѦ&= �S������H.2�d�_qk���"���.�|�����|:��b����t�Y^�������b�"�X���B�	U��)�&�V�ڎxO��Մ�m��X������A��:�ݜvQá)7�o������i2�Τ�l+�&g0�m0����jT�/9�3$�>��(���bJ�
��@�X���R���#�L�el�ȂC�Fi2'̦G5�K����x�����^f�� ��z��Q��GSK�%O�4�TP�U�ʒV~ذ�ܙM B.�>�e��Z�qϱ)'�/�Nr/���|�ز1v��h��I�?W�UL���K+�M}j\i� �1��ef���@G���$ߜ��3H��B�54��#k��2'đĜ��m�K(���7����2畃��ƥ��92춐M��>�!��m.�6�[�=�r_%����8�8|)D3�i܉�p�Ѧ����L"VJ�����z��Q]���Q��Ґ��Q���X�2{\�^�������̕V��:%פ�
�\�%4f��`�l�I���˸lā�+�т^��'�?THND�u����v:���y�`z��d����*@|�O���ػT �1bؗ�K|�#����lA]ǹ��i�,{�g7���?���$�ɴ7��?;�bwP���@�Y�����Kc"���1�+]���?�k��FT����+�$#ڜT�����	G��E-�_���@z1�.�2��{�&A��O���1�4V�`Dn�ƕ^8���2;�Z5XE��fR�Ӊk]3a�2����IU���j�V�umm��x�J'm�H"�SZ�d��f��v��hHq.::k�魀$����{�^�S�QI�R�������A��<ݎ�m�W@��pV��Wc���? ǮG�L�~1`ɻ��	
|MzxA.�+$�<�O첆/\�^3��H����^�0D,�9�UO�� 1H�z��m��@i~T6��ғ�����&�������wZ����@HG4�ZtީPQ�p#xZ��h�Х���%�Ƹ�
I��g�
T��|���6� d&\������W�
��E+�s7ڴ��/�8��AR�_k,�X UVįN=f�d����i���Yh����[��/���8$½~X1�GJ�𑢸�F"��BU0T��D�s_�֮l>�bs��q��%�w���e������*�_�X��P~0ti_U���}�m3c��(���\n���m3Q�q�Z��I�S��c(��Қ��9ܢ>�lyN`Y-7z�9�	.��=$����ĭ�oe�?���r4����;7~�Ccc��tN�ac'�[���VI�]�ܣ������g<��B.�����:��������c]�x�j���d#��%L��j�J�,�L>>���d$7e����O�̛ wךt�]���*��g���]*��|�M���Z�шiO&Z of�Xa��w�-�s����|}eVHR�RK��/��zE�>�$R�*(�Y��K.�������Qg���zQ�
#ݚ���5��bH�$�\|�!Ӝ�{64ч�G�!T��2�՝��=�oK�%��y�1M�x�@�,e�TJiQ�wk��?�"��9�P���|Du�s�,��3`N����G���k�˃ޟ��&���@�V�I�0�`��3N�ng��lv��u���-�\�c]��M���hA־�)G��x��?G�t(��3����37����r����я�.�M4��B�p2
[���:@w�E<&VcN�>ͽ�-3�NN�'���Y� ��Dc����z�Yj{|���e�&4F�`�k�[1��/zv�ycZ��^�����ߢ*�!C��x���'��k�f�,�O�p�c�K�r,�y�fo��yx׏�ތ�`z�a� ��ƿ��hS�%4b��}3:
��9'3���N������l��1�cy�ߜ�^�ٜ���?�8˥�|�{��pC޻��+�V�M4f�r�rs�������E�G��"�Vg�fh�i�'��Ԥ��\1r�F�����9i�uו����@�'��/���X9�@8�ui���;Ӥ%�.�����&.j9�����L���-5���i��<�Hz��Zr{ʠ�.�s�UҕV��Ȣ�b�ß�5L�ЙF��SLR�# �0o<�%Dķw�v�4g�i��/T�ڝE�)��D��Y�J}.�@6�G�����>��\��7��ڒ��=C@=�g�"Ġ�#����;9Tӑ�2�SD'�:C���_�8���?�C�@���.?5n):�>V/����p׶$D+פ�-��55I,QҚ��5��U%����Eۀ�e�t(YkO�\k6P��.���%�����n����L	���j�z�t�l�H�VNu�xy��H4��G���I��1��)��!T���`m��%a/O,�{Θ~�o~o^6��'��C�G�5�8����0�󢵖�ZXI�qY\dm���6=j�+������;8��X����T��0�H�� 8���y��Xri ���~����e���7y��R�F���U?DE|sq��7�0D��d�ը3*�cH
z��T�b�a�a�TV�`ă�yR��e��7GY�jb��x���mğ]�UQ^��o��/�J�M�^�˖e����8�ҍtl�E�g�ρ!!�M{��e3�F^�����)�}}�"����֓��W.8N
p��Y
�&Sš���P�׈��Ø��/��H�=2b��d�ӛ��t�F㊄�o~z��ca;6��C�5B�:=���HG�7%��Y�>.��*�V�k��/'R�M� �,�E���T9��Gߒ��dyv�3�!k ����N\,f��eL_�M	gr"�������ڞ^�H�,���<	<;�l��ʬ����t�ܙ�	����0B�K�p]����=���1ž��R��[:���:�_
o_J_��8��RigG"�����=>��q�:�]�~�����'G��MՁJ���CX$Wx��Ѡ���-���)�a�j̾�C��6jlG�e#�Yo�'nca�W|��^`MW�h�R���5x��C��,J��Eݝ�˅�~���`@�Z��=j��Oi��3�Od�� �����(PwD�XN�*�.h�o��q�o��#�=�-�wD5��eں�t���f��X����XX�/7�n#o$���-��f���Sa�+��pNl,	f�4+@�Շ>'o�˧�9=��F��`����r���?�.�vP�A�p��j^ԇғ��}�]<5M{�c����Fa��K�l�.�N���Ѭ��WV䌃�Z"{�W���9&�rZn��� ��FЏ�۶����EaUPC=���(��)v�(���9������2U�c�o���]�I��la^Q��
���÷M!aǨ:9:��+7�0TA	lt��Y�8�y��7�b�N��1��$bč�6=�đ��<�'wJ�ߝHYw_1�V�����[[k�1^�8XK?3��z����f�m&#���F����Y�-�t.ޘ��&�܃�bmlc��'<��ի�J��24M~��^�%�۬}���s��m��E�Z�bTU�C�NX����%�B�<��#0�\IR�񆏒E���E��#J�Q�	�YGY�N���~����{���pz!���Z#p���ň��Dգ�S��[��r��y��V�����w�z�W�S���m�Q�Ɉ�y8$oѣHS��l
$�a��q*у;S:v?Ŀ�Q��n5�ն0?�V\��j/"���[��j>z���;5�e~�V��yd����Q�7�tT�u�h�ȯ����uAz��18�:�Rct�M��~���#pϸu҃���f�Y���FT�����f-O�j�v
���WZ-��QRwn!>T�o��|�,D3u�����G2S��0�WXx� �<yRxA��4�zgM�"�w����0�k@z�Ö09<�>�FƁnI�	�_�VeOlZ$ 9��I�x�A���g���+�m-�x<�e��py`�%"äR!P�	�TQ?�\�
��s�-5��5k3�lYz�`���;a-�eP�F_]��]ÌZ�	<���LK/s�RH;|����v��$��Ѥ��n���³�U'���uF�� _��� �P}C��Mh�P��i��h�F���4���<�C�����!����lp�|��_T*��Q	
%Ӎ����%�p��Wq3�쿌��)O	�����T���5@��w04D95��c����2�GcGQu�S�ɛ.���f�n۟d@�3'��	M�C�1$}���:r�����i�7�����A<	ʅ��p�/y` �
 ��+�ѷ�&~.�t�ClR̨��WlS@P
;��(̛�Q�A��ħ=��V�hM�y8�j&�m6 ��~-U�"�vq_0nW�e3����v8OK���� ���^�sʀ��=�~2г-l�:)����o!C�Q��f�����=.�����5H�]�Sf	���nV(-����c4�HaQ.0�n;G����:Յ���1�㖦��Y��N��h`V�ӎ m?��|KHV�=%�:VbURc�"���E�sM��_��Ęu��N��>���x��߀��(xJ�Zd~Wu��- S^��	�Y`;����\gi�N����ZU��l�5��p�$�}�v�^���8�x��y��7`���Uv#-,x��A4�'j�ᴡ[϶����b��Pk&ߴ[�ፄ!�|�Egu}vuB��Z�|�NU0������l$�
����QB&����Ika���S�/_LBZ9K�ק֞��ql�<�'g1cjp��L�������<=�eI���N�r�9�	�n����DOL������8�'�s�ٽ����y���$�o�=WqV{��Z�l���x�C����ܤ��.7)ow�v��~�b��;��6_����bʏ��Z�OM��.-U=���3��?leAc���2g^G������V���@s�dP�	�E��+I���o�&��(X��<�ɖ��'�ĭz�/�w�zDq�co`Ήa����c.���5�zQ��e.7(�e@\P|�L�~���A�Xy��AnYP��e�8��2���j��O�YiG�u���$C�5�l��l�q$"�`���N���q�@6�݂�2�U������U5���0_M���b��?_{����l�FK��OWK�8�=�/�5sʕh��g�9�BDp�L�|D)��n�7���������S$����B
����!�W K�i����P/�d��c�$��8Pob����f��PͥVr;�V��X�s6É����I��<����2z� uq��g�I�q]�s�����IQʁP���sAQ��!�SgC_>��4���؂���3�11�࿤�Z��}��Lj�L�&#���v{3ѥ{��'��*CV'������cC�SA%U��=�Z�Xk���
̠f��q�}��O�q�ua�uj�"x�9-ES���xI�v#��4`Cː�(D����Ēa���L����4���˯Y)�m9�X�5�ǜi��M��׮`�%3��ڼ�[���!�G�O.u��8�Vh��$6"�W�w�:x��0f�\�k�����A	�yO`P�fh������ ��'kz��シF{��9{W~�裡��
o�h,��v[�S:*O�/�C���{A����
�i0{��׬<!��H,�~��%Y���%B^�N����$w�]�h��/oM�xMs7Y>?NV%��	��N� hF�M~�Ș����.��DY��Z�3p:���  ���$rҾ�x�G\��o����*8ԗ}���5�9'�b��A�����$V�R��k�	fg�0sN�: �r�{,�T��K�ME_$�uYۮ�Η}bC2 I���������,��*&���7���g
����{��^�RQ���1Q��gQ�Q��^�H��!Ɍ�����#rȟ���;$�ۦM�	N}+��;�R����S�ɦ�h�F�m���F�v^ޑ�PKĤ�Ń���a�;)�CA-����w,����^M$�{3�|�°�Y��`{̦�D�IZ��" ?k��i���p��;�'#C�H��1�B8@�������Qh��UyX$a�A�W�c������l�n�f-��(0�5r9�hh.�P�9v㆒��/��,o�yRmYܥ��U���=�U|�pBD��!(%��������9S��B9%�2�7�]v\J �#;���@�Z]�#=����MR�Hܰ3�%�)�N��E����'@��j3e1�Jۡ\�U(4,�c �}ܭ(p�&�a��Ŷ�˞q	�%8�x�S���1i<�E�|�ǜ�L��G��up�r�pQuy>Q��2��c�ZH�d�X�����2�\�j��5O)��9�������ҙ���:�"[�"Iψ
�������X�)��N�Ҩ=�%���j���+~�#��R�c�TE��\�h�N$Z4�o'l�Yn.�������]���Ky$b�C���{WC���%c$�`���̸�Ê]��Պ.��6�Rײ�����AF�$�a�+"��	�/�0�
�]�K�c�0 uN��c�,B�y���dF61�O���F���5Aoe�9oTx!��+�F/ڸ~�52JꧩG��t-~8�q|�<��s��t^n9&_�BP�E��̍�T�͐��?y��K�FR��������M�'	w��UW@���p[=���B�[�9%�O�w���2��x��eM)�V�֩�����o�5qk�aL��C�F�P����%�J��(W�T6��������zwW��?^a����"�@����F^i�U�'y��RM�Y�58���x��>��v�X# 
�����^qAR-�����MKP�|9+�����nw�LD>�AH��i�Uk��4���+OO�_Y��S���!P!���p����ắy�S����K��s6�`�K�)R��,�~b7Qg�"�b��t�"�����2�?SZ���E#�?�A!�7Q1G^�G�=W���)��'��;��������^����j�e`%Z��]������~���_0�[$+�<i}K[b������m� �O�|r}��|��q玛^;���6�I�!��>�ǌ-���Y|����Һ�jȱ��o�d֑���B���b��o����ŷ$�ѧ=��"]��oX%���*wdЏ(i9�R�@��ss��:�]�3�$7�*f��w�M��ȕw�ཉ���y
���5�|M�p���d�\�僚�WnS�����Գ�[s�)��f��xpn��
��h0'����l���a+:O�Np: ���d��g��������W��Z�E��#�:eY|�19��(�i.��ᙍ�[@b4�;�q�Xs�(Yo�p�+H=�~W�ƯI��Y�"��B̡r�� %��d�v;&}��}�Iz�� ?0('8т,���?>B<?>�/�
KB��w�d�n5�A^d��!���{8���p � �_Ԁ��bh�&׳4P��̮j��.�HA�хQ =uԩ���}%k�vg\����X7�B��-�P �g#�ծ�n�֭N��w є�j��;��zꋙ��'�b�����H�+�zR]�3�?���bHN��4�J咴���UH�}$�7^7�i������|���~��B�ߩ��k��|� �1�@�[IP��R�3#�ц8�/A���#C��Jb|���R�g� �Q�W���a����!���e.�H_^��S_�o���c��>��e��~S��m�9J��%s.�0p ��J�xk�OB9DyQ�F?c:�87U�6p�YYg�������d3 �Ϙ�A��a�����W�l[m]�(r�)c4I�u�T����1ڂ�'���D��0g?����'��Qm�"<l?����%𷼑��J��װ]�g����q�ҟ���0 1D�.=�ݑ'��	��9e���B��o�mbe~R5l�Ѷ|R��'ʣ���̭�+�	�!�4��t�‪u{l���K��:�"�xE�Q2�'	��ݩ���S'�ɏ��8��c��m���_j����1�Ń>�ZY��E����^���J#ĈW��2��
�OK�/7�$6�d�C��l�b�v�*�����WxfP�I�@�Brm1����x$2�:�@N����Y6>G��[�{R�� ���VN'��#.N�M����;��j���Y��%[Y 6�*Ѧ���o\�B��o�o�k�Q�#��љ�		�n����*��>����_�;����7y��C���X���/'ms2a���-� O��GL�%Fa�ce����7⷗�U��X�7���>����M�(0� �(���W�=ۀ H*�[@�->�H��WZ���Q�Fx��L6T��l�H�g�¦6OUޑ8��3#"BN�zZ��gq��.S�X��Z���ψ�W67k��2��D���OML�gV�����>����dqa���#�5�w��ŋ��J���eX5^iDՕ-r҅�@?��|%�b��>~������ټ7�J�d�:���!&�����Jh����#������<���J�;~7]$ �zd`|��BI!-�qkR��E��U��mn���/ɨP�Ǹ��������0-�l�����\����O=�df��'t���£�b|�r��s��� f0�)-��# 7�Ϣ�t���&.��nF�
�\�ZHIHpZ��~3�� (u����"��`��v�m^7��c�*=���Qys�m��]�ѝ(4��R�W��ݱޝ�2ە} A��
R�>�y�j�����=$����c�=±�� �٨��+4�b�-�6�0�v9�2�$��י��E,@5Z1���p����,����6*Zt"v���ek���6k� $���TC�#�j2����!z�'���P��a$ �,o|=��u�~��5@�/���>7��Q! t���NhL�Ow$��:�������}`��( j���<4���y��zĻ,�_�!j��U�]Z��}|\��P�>��dLӰ,&��3.Ep�J[.-?�|�e6^�Ů�
�3y� �b����7��{�*߯��U�5}%�g/��[��-�"9�r��w�fR~_��+#8o,++7L�d1��*.�2�C�>!Lb����Y����1��Ϊ@J � ex��t�|%�W@Od0S ��i��J���-��T?.~)�v�T7H�kQ>�]?�l�W����4�k��� �X����ԫ8�[�����)��Ty��V��-��~��g҂�z.h�qӠ��[�Ls���}�g*���Dm�9p3�W5��%>�F��JW�&+�S�L��O�a�d��[�N�Y�P�@�c��#@�`�H�{�2f"t�?�X	�D!zw�i���t�<�gM���c$���0�K�����P�R�/[id�W�,���u^�I۷��Yvc�5m��ټ��opb���#�2�Lns��q>�l#�$���u���0=O4��q�KH~��/�o��bz�7�x�\0�&mQ_m{�!�Y�*,T�R��6TQe�@6LH�����~k� e�2B�N~(y�f��td�?��'9��}�D�E���{Ă̽�r�=�Z����Rcb�.ú"���Kȥ�$�5|��gCE�$n ��e��푖�iH�3���@��
s���{�� �I�`.���'Q��1�pNa\��H��aҕ���Ri�����%Rn 1轸�.��.2��H7��7+YA�C)4�˙�d��ʅtn��(�۹x��C��U��Ě��A���C�p~g�*�Ҫ:^!���:b��V�y ֤��i�1cH�A����M��d��p�Ĉ�b��!�,;����|�!���z+F��,�7<��U�u�t;D,#�	#�����Ӟ^(>nl�	9����E��6��ͥ�8INʌ�����iGۤ��코 @r�����/��J%�2���Wj���v]Յ�P�w���nT9������4�bM�#�5�xb��N)��'�)�����I���B��6L��=��/<e�57V�Rg��CwS/�C��"f���3�`�ԬVJ�e=���u�uH��OЫ�"������`gEr��8�T���r��J���)��wZp�E��@M���6�K��;J�������p����ie��F-���3B��c9��2��&��ٟ�����	�ヷ�� o����Y2��%Ĭ��3�u���桥��
�D���	#���2	,f��{]S��v#����F� ���5�&�n����������Qgn�ִd��� !���'�]a�&�v>z���h�y��Rkp`ݔ�[�\�o�N�lT��
d�T2�a���D'2(�p�P�w'����C���8BWf���޺(6m��*1�%�[��z�f�:[�*��!�d�̏���VE�tL �sS!j�����
ى������/�e�hp+�V�X���la�\@���<����_��7���bБ�>�:�(,�g�d����Y_�;ݞ[���.
��y�gUe�Z;�+�$��S٩/���=��R ���H''B�Z��b$�	��p�v7��UK������^ȸwau	����H�p�I����D�q�.&��.=�H-+e�����6��:�W�a
M�{�q��PM.p�R}�Y�k����G�7r�[U�Sa�w�!m����x�=v��}\ȹsA�u"U��Yfu�t�ꀃ3Gm�*Kz�Z������9��n t�:����4)����h��{���)1t������w��9�~��}ђ�0`��xwu���u|I���\:�i����(�n���,�獥�4B����R��A�*f��I��,}r�̷9d�HB1v����|�0D*�Fܴ��� F��/m�qc-,=vl�aQ��MZ�����ۤ�i�ϰ�)�b����Y�:�O�;�l�Ѫ?���,|��婵���Q(^&�OQ{Pv=��^f��ja����9�1Q�]��)�[Ac��4���ٽ�1NH˧|��>S��o�g`�|Z5y1�2)������q���a?ǆ14�Q:�г���v�m�@�J%��凷�bF��%-���[������;�����R3c��?j��ݍ����G�Ǐ��4��
���29��=S���|�����#(M���g�2��PD��6lE4Z5�5��%�]�l#���A][�ؚO��3�c�gER)�B�}z:�$��Z�`݅Ŝ�F�m�iSw��Z�ܐ�*�!����$ܸ.x��Q��7�+m��]$����c��I�"��U�<��pE>��F��t�����9�%�wp\cֈ�޽c��ecK+���w ��;f\s���_����A�P��I?ޗ3����n/�1��M�~_~�O��v��S�d$�E8HU�_>cKv�l�1?�t��u�	>^�6VQX�p�^����y�V��^��c�s�@���D�P�OA0J^V�t��荡�C����v�OH���
�gO%u�}G��?cߋY�G��0��(�hG��[��сn`: �������ˬ��<+A�׭F�	�y"
<	�Vyz����;�Cf2� mB����rm,�FZk&�{���1�#� l�!�����
2�����/�r��	���<��	�+bT$�M��c����i�("�� ����M����`�7G���:A	��"�y�qr.$Sx������+Ɖ�u���H��`�"b0���Ό�}���R�������zvڡ���5]��#�*X�ޖ1%��J�Y��M�����V�`�D~�f��M�y�:�GGo����&��p��7(���B�*�!�I|�z�LM���e?����]Igp]'1���)�Լ��}!l�6d�+o	�`���A'LR�5��g�;9Y�Yi>M�l���)�B���H]��C�1_.�	��`�a���?d��{����W	��Y�B�����&ǝ������	�m����mee ߈d��)Ϛc?W�u�+��D�5ޅ�ܜgڐ�L�JCͷ�vX����F��t�eh������r�!��e��:V�5L�� �СL@�� �R�!��A�x�ё"=qԴ����֟'�t�⻗}zP�10��P�r<��,�.��[A3ˠw~��#��(�k[b]�l�q�Θ2�g��Pu�x$ܑс����|8{��A�E�����9E��JU�&����=�vP��/�:(�4��ڸ��uq���l�O��W�%�:���WT����ܦ�'�g@~� ���h�)�˶Z	�bى� cC�Ah\e���%e�,�4�8��y��;��?2Q]�+8]�;*zo�$�c�&�I���?O�lX������E_�[��Wy�f��3��a��@�-�[C�@���Ǩ�'Z�kT�"�I� �~�=�@�ʊCz�H��7�U��#`Q�4�����2ۇ�Y<���(�S*������q�dB�|d%��?1ں¿�)E,?VF��7��t|������8ew����x>���9���o)��60��RQ�y�w5y���҅^cn�!rjK�Q����<�Z��t�D��<rg_���g�}�r�� &�����χ�<��-�4��R���C�׃�G�M9�}+l��(���.��
E±�~�"n��uM�o�_�򾘫��(CR���2��ȯL'{���_��.ܤ)Yʁ�I,�S�h�KD�a�9M�� ��敜x���jO�Y�,�@S#9���L�=\M�X���zO����j&�ٵ[m�޶5��z
���dn��$��d�jA�|T󐊉��]��]������v�j����m��	V[^69Y&�q[�mV㐱;�\��dͬ9mtV����f�R�q��8��I��N_�����>�������U��H�����፷&��[�Xo��6�� ~4������^Z�|����m	�L`	�) oQ߲LW.A�?��R���M����nѻI:wM�/�u�J��ػ�1 യ�h� �"�y��w@[{�C0����؀��ar Ra�AO���_��f�#��4U����MN�D�2'��Nb��y�^8Ք����J�����(v&i4/���3r4�� �����^�Z��ja��G�ST����c�ޕ m1$?=�	�Σ�\�K8a`���.H<:�w����v��Ű�]��Q%:mJW��k
/������d⤡��Աoת��a0W�y�0�bB-8ɥd_z�[�׺]���l�ʚB�F��(�ˈp��eueQ�&X9���tE]���r�}Dp���g�f�`�;5;�Ŝ��Z��@uB��C|5!�'e2%?�VH���ʆs]�I��[�{�j<�=u�b���5��sۢ�e�VVu��{%�r�Ro�U� pa��[�3r]+����d��Tt�q8���V�h�ör4��J���D²c2M���j��FU�K9��>ω����0b8'��s^m;4�6�Ȯ!�X��T�k�*)w�?�tO^���*"��! �ߩǋ6��/[�J����1DL����<VDQ�bw��[|��`��-n�lXfݬ-�ʙ�]�r��N��^��� �|PQJ;��Lc�������K�鞧�T�%�⵷[��G]�����QNc���m>�81��ǘ�������u�?���g[���W�������ah�֍�]�����ͻ&[�u}U�����m��y��bCJ�c��������a�`PF��%�!|)��{<`վ��Rk6�m�i�
O����qhO��!��MqW)��ӻ�V$;j��{5�fJ��.���bǙL�H���2��x	U �H�`3�|����  բ���u�� mPr�}�4��bږ����`��s���� ��k�N�����2?9�I��?���@��i[�ˊ�3�����6Q��Z|郂�8i��5��a�I���U�*�&گ���M���I^�����Qfh)zt�E�]������R�.�HvEk����q�|�SY[}�^���*:ݾ0 �+�V�n@w"
R���oc]a�������r]^�e��\�<$�Ƹ�`��Ha�����g��%�	kX�E��s,xP������"��ǘz��V�ʌ�s���������o�t��P���0)�dRl�h���c��Ɍ�Ȋ�%��JI�y�-��5���t�>|P�����W�z'#u�2���s��G�5��LV&��!�)i��|�0�����Ft���V�ܥ])9R2�Yp�7Wa5�e����s��Oчl��U7,c�/w�nm�+�� �7�=�e���Na{�O�78ۊ �U�,�S��;T��E*�	ŃJ����'�V��hi�7�崅�1��Kf�;��F�XF'o�2�6*z�lͭp��;X��w� �(J�Q~��j?��>���0c�=�l�yeQ��~�ok�� ��x�+�rdpq	H�_�O�� :�5��r?,���b*�I�4���Z6��:b7���v
�;v����H����kG�GO�LV1zo��؟������ݿ��
@��>�:���>8vIqP��( �����4���x6�:K�[L'�,�h�ᆐ)�l��{���_�#沤���d�\���xQ�?*����$ �L
O��T��+)B���ώ���w�u?��hn����l���&м�.T���$sz�P`
�S�`:�T `���
V�p��"�)�� �b���vp����1Ht��5��sܥq�b��Ve���S������:�!�=ֱۋP����-���V���衶�6���C�z[����c�+�m��&>$�E��dѸ�Z��r�0(-�>�Az���M��M�Jeƚ�o��W��ֱ%��� \A�FEg
D����$Y�*�S��R̮�ÝO-{K(��)���9�$;���_c��ꗵ���I�u������KԲ��#��Li���PB'Շ��1@�7e:v��$��4��"�ka�W_	�+EAJ.S����֮e�ƶ��V�ȥL��N���s`�R$� �m.�������/�7�i�|��Y��k#�ҧ�jf�e�#�K��u�Gh����>�GN�7��f͖H�ʘ�ìg{0�~��HuR���̧�|bU���
����ԉ����QG�}��(�h�/'�+Ul~`1��H^]��<J���ur7�>��ʎM�8+�B�PI�%��i�b̂� V�1�bC�i�Bp<���	:��.iF~ X�|o���-�Y\Q�Ѯ��k�
�JE7ɟ�����^T�0��~ź�JG+�D^�1v^:8΀J��C5h�������sO<����p��'��RD)uW�x#�Ʀ��_�x#@��[��7���<*��KQ�ky{�}�Gc�r8�#�� ��D���@�)ȷ��|m�l�nb�Go7��R����IV��:ƺ�m
�^�˞|XCr\ŷ]��������V����|����H�V��|$�x� #ƫ0��aW��2��K����q#��Y���n\�A����2�?|�J-���˾�t��"vG�vd��"��{_'@��Q�5���h�*��:~f  ��(�}�D@Ix���97�<��}ʵ�q�D�ٛ�fL 5n�D�y���T��<�+���y�|&�%3a�c�FA܀��'dB�1��0��!%=H�Z�'���ŋG6Ɏ�����
3�~�8�o(ց͖��;�<�(�#n-�c��f9kt�����0�*|XX"k��К]T��UGd�-� �:�w��ܭ���\"��F�<�|�}J�u��<�У�����:�������	V*s35��u;�p�QF������&~����r>�\�k��R�>��Q����V�y�?@��~��dl��&��7�[���V���u��$uh���2����ɫ6N0��,��Ԃ8�nBj�Ym���g���
@v��?������	6e��1o�V8�8/%��r/����8h�Փ�qgI��K���?�z�-�7謷"Do�v��)Z�H�u��f�Yiuh���g&�r��h� ��5�;���HI_�1��C�ˌ�n�k��wm�� y��
x����1L%`~��a� x���~k]|A_�k �M���f�*�*s�WZS�%�^^��Gg{�r��T
UE_K�_����������U����2?��Ӵ�?o�DA���WT�n�xA(�Trc	t�cWյ��n��'�̆6�P':��k
�s�oB1�J�Y���$�B�=&
���I�̷��T�T��S�R��M�,r"��aq��Z��d��2T��4J'ZM��� �|bN�ǵT�����U�-4��_Wv��I���_|щ��t�p'o��\�5#���5�xvر'��h�:��ۏD��V�z��Bu ��PX���޸�J��1-����/�{�R{�,��F�.�mQ8�h&��\�S/�&ld���N6��{�E$��i��A��sY���V:�ٜ<��jB�A#Vi0z=�]�q��arU1Vb�M�3�
��`�3�W����Qi
Ց\0��
}�������*Н`��=͙ �_��&c���ca��~�c<v��d%@�k�ᖦK��M���t���t����aV�\߫�1������x�f��h.���4�_�GML���X$���0T`u��)��d����vf��	7�	AYp��j��؊��Oy�ˬ;H�����㸳Oum��5�����26���lݣ-�O1�}�7�Ä �V�FfXiV ���{07�$
.�Ls��C�|��*���w]}�@�3̢9�F]$/�i���9��Hs�����8حʒ��5 Z�p	�0���%�uf�T"Op�Y�%�p9���io(�d�a!��I����̐��x�g�6��PN�~��%��\t�K>�e��HN����l� �T���"� R�l����G䏘'z��(@l�JS�70,u���tF�MK��O��&6�DY��x�����y����
q o�-�w�a��魾���\�04�}�ì��#]�z��r����6@�ۭx{
�������5�]=xC�gg��������u�+r-A��w��°�=�E|y?7J��c[���U?��u5��-(�<�^J����3�[�Gu�q��C�� }\c����`�H�
}����3`:tY�-�g��K�a$��7��!0�#s��Z�L�	�١����Kz4��~�"�1�YЯݽ\֍�1�k�<��q)�j�x�\�z�',�x� ��Q�t_L����nyj!c��jh5�xW݀�&��Cn&LA�卉�6�[9�CBG?9�v�G]��%�b0���w�����p�R����~��w��R�E�L�%�!�O��	,�/�'���r����<g2)��X1,u�p}���r{����`���s<��ސq�;����	��Hٶ�q�뭥1�X���f���L���-E��ЀΗA�R�#�d�HB�%�͎3���˥4K/x�	� (�[S�ni+�>~[kn �HM���-�GH= �~ɦi���-5���������x��OM�^�������[}�aϋXJt�A��C�o#d��<�"�@�Q� ��iu6�&k�f~%�C�!;�oqq
��T�F}��0=al,�aQp픁.ʐ+�g��<�Y`�5��>�C�v���}jT�ȋ�`�����3~F=/E�5�z�C�Uo9�< W5.-��>�8�-���΋���z�ir\�AP�u`-�����M�X��l�=����꯹�\�r��i��(�;M�������T��Ok# �ƺ<�!#߫͐��f�/ĭ�?�^��_;F��?i�^<'G(�|�$��H�����,9�e��v'�~MXr�f1á2����0A
�æ���v�~�#}:�~�V�]�<�s��ǌ�PfrH��� �1� �
���ۋ&�'/j�l@�L����q�:O~���$@�������j��쬹v������ ̲çI�1�6X�:R|�B	.N�G�����(U��9�,pر������$T�[��LB�2�m������ZE��r@�+��L�¼l�Җ�b`l�}�Zu�x�+׀{��&HizᚹI���m�X+bwX�ȿ]ȉg�
��Y�G���X@�dzG����b�<�[ȌR����e�sa���]%������	&��>��!a��"��{���FaRK� ����W��n]{��_���M��C
��#�����M�Y�x3����_��p,����e�����?�ag �pJ�	j߂�%vU!��өB/�v�?�قՏ��,�p���VOF�50!7�b����1��V4ZW�>R�퍦SEf�#j�AՒ��	�ߝ�?���b��MS8.�pb�/<7�˓ܺ�����M݈����j�<T_��m.���K�4J1b܋oJڊ�����9�؉bH��Ѩ�k�g�n�}�����7���_s*݃I��I6뗼ߨ{DY�C  H��}�l�eA�dW����;`& 8��i�F�����˴J��i�4��*W�=��4�WT��
S0��_��A��x�`�'�w�\�.襅wk����s�!��YF� ��{��Ǖ�d��?U���]��Z���.8@G��.�����F�do��:3�Ǆ^�;�׎�iέ���dm��o���l�F�߷O����tY�lQZl>_���W��;k�LLڣ�.ۻAߺ��>�\Ff|���;ّKx)Ф�P1��и*��+�1���Ӷ(<��k׺
B�M������x�iN�O��KM�\%B�jْf�fri�PXE���d��y��:/� Lӥ�k@t�;�g������)�,*-�r���sӟ��9���蘝ۧ1�����ģ��Yϡyv�D��9���qD���O�M�&L!�`D�����d��ۙ����e�.�xR��p_�w�x�|H��~��c��m�>7u!�҈	|[)G(҆�̧7bu�C�VRH���bd9���LR5���� �S����n�
���$�5�Ğ���YU�0��q���W�)���K3a�B���N=Js����a3e��+�uLP� *���c�[��t��Uf	��q����ןD�@��Y8���5?�1���,������wL�K��T�����*G8�w>4�fW�
BTRB[k��.�[8�+�@tU�ސ,5�����@[�h�FB����r�b���K����xb�,N��j���f���kuE��q�)YDZ-�<�zz��A��mŧ�A �Pd��(��$8��+,桱�̵�#	Y�$�:\���k��B�WH�]��m�S+K�|dF�_����#���u�;@wnV��3ȝ6�^�O23�hDohSϮ���,XY�xl/n��;�-d�V��J?ĨMF��9]�c��n<͔V�V��tL��҇�G��<�`�5�)�|��%ޱ:Zޚ�U��ң�"�'�	Y�?��(��� �!���VSM��I����,���wB���p�e�����4�0�5l����C�Kna�<^x"""�d�o{8V6n��1�[�õ� ���������r�*os%�ǿ:'�<]t��K[�Y�w�g[I�OK����ý�9�fp���pЩ��W��wO�'�b7�q[�ԥX��٩>�L304<�|���kCpIs�)��1;�Yjj�w���K� z:�:=�S�aT�wˬ�~���M�+HyJ����7>�$�Ӛ��ù��_dLv �땹 �W���.��=��<����8� �HM�$�$��'�U�M̂q�eQiU���8f�Jg54&$HܷB����H�f\�[�Rr�p��au��B��� (���bֿ��@5\7eT �g��OL��L���2�s��q(9ьxv��Ι�KuMA94�E�6������5�2���WU�;���#{�i"���AÚ�甘���<������D��
��Í�
�'�I�'y%?$�j��.?Q}@6����*�vv"����U��O������B�"��$���� �;�$%��ZW�%5���/xs%L��Xet9���%��1F[Q�6�Q���NOPT����Tq��UH�RDC���1�x�	w��"pL:]ԇ;���F���N/���=$���46o?T��@�o/��諤m���J��s�AWY�!��a�R�>���� 0�b�MK��7��T�p��TAj*��J���F����5d��R���czKD��$Dp�xk��>W�H'���#/3x�q�C������u8���}� ��'��݄��R�OX�6�S0;\a�)���Q{��Бja\�ֶ|�.��;�׆���	0��!�T�_#���k*�7���q�-���"g��ZX��fc�I� ����������fp���c�c�Fg�,z�����2?��゚����j'2l`�0kK����"�Z�fY5��|B0��)���b蚝��g��R��-����O�Ј1CUG�w�f�M�@:�("��azLIB�Y#U٠M�\w�o�գ����m����WH��SL�!Zcq(���0�g8$&3���\�J豃�%�Í����
q�pF���p8�PX�_�:�/'��#)��4�c�!���Tol&I3E����f$���`�C�)I�Ϙ�/���4�8��������g�z�gK��C�t�r�_��b9�]`�O+%آf��,o1��].kak2SF�YC���44,e�hӁ׫g�<�@]���SoI0���Z�<�M	ಿ���;�͘���S��)?H3:W�/��c�0@b��_�R��XL*͏g��\�����������/H*�'�<B�Gѡ��p�}`�0�0D��G^g��X����]~+v$W$��N|�hMĮ��"~��\�7�Ybc{�x�.l�� c2��m��uS^��>�j<�#L/�B���&W:A ��3^˥Ϥf���K}#_$%	4���P1݃]8�� �R������j�ة��=����cF���
�bU�r�Y����n2��]�}��-��@�%��J}���gAc��l��$�8�
?��JH9�}3:|��#��%lI(v�>ZR�]hNX�Q��8-�S�ѿ��0���y�Ahq"FP�:ǣ������?���G4q��V�{�(�:�����lOk���b
�B�2����sv���~��-���z��(����YENN���y�͗��sԼ��B��Jr�90� ��P$'�|ڴm���c��ʓ�Hu2 �g�����Ѐ?�U�������(��`�y[�Q�?b�e�.V����!��k��-T%P�s��q��BV�����̀�Q�Ö�uq��a�M��|+�⓶�x\��:��N&�P��x�Ƙ�A��9�qE�\,���n��*����v��l^�]z���w!�=��O�|��?{b)^�P�>\iXeE�%#��5�.�Ҷ�p�@� �ͯ���I���zY� �8W{��@���v�a�\" �������OlY�	<�>�������^Ů�Q!6s��"Y>�yD2;_@;1^bE�:Uq�r����d����=������n�+��%H���~<�Nة��3�X��ZH�M���u&��f�i�����,��'<k!�q���|���f�濉��5�2�	BHY�7�����g*]��-w�z^.��C�oY�q�������p���D�9��G������Q�E$��O�j�n0�3,?���ō�����O�)}�t�;'!�&��i�WT���8�M���v����/�̖�I)��h�@۶��p��p�HXʔ�J 3S�����ˣ�Zu�ֿ
���3ȯ��1좧/3�~O�0��l�V��}l��s ���i�1D� ����cC��v������\0�5�1GRt\�
N��0�=�M�G���	�9n��L�����L��30����qS0
�y���ց"_�����ȾxZT�Ŋ����;�!�өe�	�J�Gq�J_-�*�ˬV���i��I��ߌ�/-�x��!�ӊ�x����_t��2b~I��vQʊ�Hx��h�.��h��ub''��4��۴������L�:G��5��,`�7��`JV4��t6/��x�pm؋t��_.l*�3�c���Q"ף��6O�|[�Mo��l�r�I?�DYoT��ϙV"���"�/�d�@�,V���d(wɯ|l�! �.�o����x`6�Z���G�ڃ�[t���t�./pMеn�2��$�v�|/���lʌY��ܡ���"���L\@��Ú�����X�	 3�GQ߇��U������[Z=u��fd���#=��Ք�N�S�q�4��l;�Í��rF�����IJsR�Ĉ0p�Ĥ�.���)
�1orw�-��ʺ�kE���$���8fe���6���:&�}��XC�� l�v���2�HE��tf���Bik�F�
������%f/`�8��D�oFlș.1�|���S[���t�ˢ^�����y��H�mx���]�-Zx�r���Q5`��i�|UV_>��|��������f@/u'(Xa2D�RW�ǽ�EUv)S�"/�I�ʨ7_�Kc�}"F�B�&�)t�+.��bU=l;�G]��Z����
������#�b��������E� �JӸ�u�P��$��)��dmE�Rɍk�ޑp���2TaRO����6z���V�n�B�����b��P7�5ctS �����o����*������u����'�r����ذ�8!I��E|�m�]���@��n�q2~����3�&FB�W썕��V�{D<=��r*d�VI{u5#�I����v0KCI�J9\�Ѐ�0����2�@'F��$�&G��S,���5pU	
��1��o�ny4+����&p!G�Ot�E
�J`ы�k�tZ�j�^qf��LІ����ܗt(Oc�e��B��\�	V�Bwqd"�3��I�������BàV|d��O�H��nq�pQ�@���-��q���R뵨�;�!��JUO�6a�<�|�o��_j*D�]�s��f|p��ߺ�!�b�p�-��2.7�hg�����{����3�*���Գ�x�����	/^�"m*��s����������`��?���0�\J���!�����11A:�4�"e/�N}A�=�A��lS��j�C�^�S��y�A5��XcUAw��|�3q"HwLO$����de���9ꞷN�M�zL��(/��u��P��U�M_�"��I�(��?�p|H=���r�p?��`v`��ُ�;�ῥ�I�7�h# DU��������9[��zХ~�'�wι�c�����#=�����?��51�Ͳ��q�ݱ�dm,S=T�ڛf7Y�oN�����σ�S=0��]�ځ�P��2�I����Y�R�� MR	fNA>7���Up8�"�Q���+q!ñ�P��ve6�`8u��Ջ��ע�	Ԯ�{���wC���1�A��V��s~�F3?Ob�;"�x��@h��Ư�_�o.��鋨�G+ug�±���Yz��^TLB��E��'q.��b��t�h ϱ���@|VܣQ������B���t�ec��)�y���.��?>p�l���!ϒ��/�f�0;�4�:u��d��_g��,�T�w�)���	�n�!�RUMO���5�s��T�@3���\(�� ')�ÿo\���J5��et�MW��r����R���T��03�qqЅy���X��JV���;��}?ɂ�e�����5���R�z�K�Uj:p�|���(�|t�Y�xX�N�]��ܩ^��b�f�P�]�֐��+�8�,���Y9*c⸗��LJ�uv↦(�B{&]�1�q~��s�7�\��gl9�<iy���([�bn�!���� �f���)�Q`�!��.�5�$�z����x4�!2Z���*Y�&�d��e����-��)�����{�X��i>��}F�p�vo�p�E�Ĵy�Y�K�����М:�%j]z��kT�x#}�hv��[�и����"��h�)i�5��������g�V��;����C�s����&���{�Pp/�ܻF�q���m����a�jݓg�O�9Q`[��"���f��LZ�u�}�_o���X�^���H��ֽ���Y��L����Z,].k����&C���:���UC�ˢ��kR���/U�Ie'�w=�C��&���m�؂FV9���Lm�g�j�!Մ�����]KZ��d\��R����|�.�����qm�k)E�Ȗ)�-������w" ����O�pjgL�AJ�*P��M��ꩀ�_չ�6;�?��\H�&����Z>�[��B='�/�p���
�����y1�>�{���RrKٗ`�F���X�9LI�S-(Aݨ��5�j}��Cy�h���ӑ]F<�N"��wC��H�9�d�����x�NH!JT���G�虳C��MX�`�!��$�� ]���2�wꓠ���Qb�
M��@,Z;iO��$�N��v���		�������v1o(l�ş���y��d�jY&Q�;0��ӥ71��\��CN�e}U�l��[�N��;��e������+��>�'�<J�G�4S�������y�� ��L7�6�~*��0(�d:d������V�1�G7��������EJ8Ke�4������H
��P��L�uO���b؝%���}:���7���lx�S����x0�$_�c	�������)m+���m�u��C@���!O��)��	XavI8�sp������woCf�yZcL��\�
&��v�����7ڐ�FU�Ҷ�S�5f޺��)��,�"�B&��Rf,?������,]��̀/$aM��@�qt/j�1O��/��yΌ�	Fp�O�{z�L.ԪA��j�����~2ҋ�j�Sj-�2����&4{��x�q�Q�$D~˩a�]ҿQٛ��g��G�/M*��d=�{GY7��8n�Ǽ���]�bu' �g�F�0�CLd%�A�����nз�Ь��5�`A<�c�TKA�Q3�AjD��ۺ�#���VQ�m�@���9��4y�[��|�m�~��S.��a�T��
��X^����>�2b���nBe� �Q�r���A��Z����Z����i�a��7��I� �5 ֬x<	ќ�^�Q�1o����\̆n6�:˧�f�7T�Xg���e�B�7������a'H�R6@�z�Y�v���`0`�KA�!l�����!�.z�&O�Γ��R�RA�q�-Y�qK�!���gĔ��j�xqC1�|� ���A����`X�&�@�:�݀3�y���s�%B��A&��N��l�+2�׀�CF�s����Hq���[��A�%����I�%ex����5"tI>/�[�*Тu���0r��0r�|�7-$�ԙ��SKFR�r�8EC=b��H5�pנT���{�!΅K9�Q0y$��J�JV�t����J�<��Č�n�	]��4̽��~�����O����}	/fS�h��|��:�;�HpЯ۳	�%U�ohS��2���W�G�Q(��Ě��f�#��(yo�\�TgA1�BQ]�	l9�ZLV��)iu�$X��F4d��T
 ������~Ǝ �R�xw0s$�E�����ś��
H�	�~,��u#]X�e�q���� ���z��_bd�[N�-Y��r:Ͱ������K&��b���y�1�WM���6��o�����- Y7�c������_$�J3���w
K���H�q~�bܻ!�TT�T�4����>Y�:W��|�@Q�X��gXo���̀B���'R�VM +��*��8*�5'�e��lت^a5=nׂ������5�'��J���yñ��	���:������v����I��+E�����>�U���Y�����^l$�U(�=����F��dRḱ�g�3��A�R\\<� 
�4�luu�"y2�@c�L:�K�t\z�=q(b�0ֽ;�#+H�IׁA�%�Syʳ	�H��
~�0��I�a�ּ�4����>������6�
�E��Oe�<�v���d:��(��[şI'd%�
�����Q/'J����4�Ww��U��Ԫ��@٠::`��F�@�%�n��Cs��;�Ahˀ�� ��_�C�5e�HZy@��y(!)M�`Vtnɂ���sнg�{�En���S}Ï� �zG��{6Qv����>0�l|0���
.�o���߬k�H�ޝ�Г���g���F�Y��1Tj�4�q���-�����s�xI$�W���z8UE�j�t��I4hkN�X EGl"�OC2d�Fд!j�#�K� X*:u�ґ<�~�1[F�K��a!Vґi:t�T�LzAfd߀P^.({�
�^�g����y��)xܲ����3���Pt��yD��)��s6�@�q�׾���C����%��2(T
I��Y�\|֫9#��>�Wƙ��U���'K��-&�[&���[�br���(�[� �xڡyA��N5��,9��{��q��E*�1�Hn����Dĉ�8�O�A�u����:�@_�o����"luKd�F�6` �O�O���L)e�U&���
.6��Ph���kh�\��*�5`���G/>Cn�}ř���_|q(?�2�'������>��-z�P�Ii�9\n�/�q�P�g�yd��\�"V~�9y:i�)�Vs�Yz�!	>6�=ka���2�⣈v3^B�WK�4�JV�N�n_���)�/P��+�T�>x[C��H�omFb9��jaݖ�@�(�˦:C�ѭ��i^���{@c��� p_D�	��ɖ��@zE�G������^ ��oahs��>q��X�����G�kY�$���$��ۆ5����9���5��5[���M��������Y�F�mP��'B]Q�o���ϵ��B�E|è���L4�����4��.��K������\���S���O^���D��_�/�k��T75e_"��YᏯ�d���f�����%�.�&�}�x���/(��P�e�`K�s���{7$4�7��Z��<j�9<MD0J�8�^��&%i��u_^�,�:t��XL�jT�I�ˉ�Ceh�B�`le\� Ҍ��Ь{!|�|�j6�_y�y!(PL�=^>Z+.Pb�Z
���k��Ɓ�;�K���܂����c ��ɗ,T��L�uf[j���Y�0����Ng��ʴb"{��
<��V��ns4��;��;�F8v2�=^�b��eO�X��Ŷ4�i�GJ�2��6�щ���J̮��=�<3s�&�w��Q�����Fqm�CN|�H3CeQ�r�>>Ip��Ig�c�/��o��
Fs����K%d��RGZ�=�%��ć�h�҂@y(!dt��� N��@>��u-��aP�j6JG`Z�[Ҩ`0S����{�|-����X����y=�&��V�,!Q�A�ƾ2��3H���L](&�� �%`�F�5/9Y�Ɔ�݃� ��(ܼ��\�8v-c�44��ǍTe4y�!�m5�a�ʉn:XV~8g��T�1�{��-h5�V�؋N���,�pԧy��%�v��Q��b���.a�'n�*h��(ú�;]^ԪQ���K�3��0�'J�噥;,��l�.�||ݥ�el�CQ`�s9?�쇂դ7{��b��;���-�غ� �mˈ8a=Eh9�	�IY|Ϳ����8qh����J��V�"}�55WyEu�FX1j���H�:�)a�>	Ewf�g�B��w�Nh��H��$S��GC��o���L*���y�^&{��H�C� >��(5���X�-�G��6M�;�t�4����ZV��T	����q'Dnٲ��k|
���s��@Cc?i��_#'6�9�Q�gK����_ݜzr�a�O|��p �q�]�bT��$(��+������	֞I�|럞l�X�{G!)�0t��^�jl��ʡC�h/���Uc�u� ԩ��o�@ /-���_wk'�FMơ��,N��]Q��"�I�6HFL�<��I�.&��o��}��Y����K����
�E�_��Z��������p���GΔ.��<����|���+;z(��k�Gb��b���7u���E��S��vϻ}�$-2o�Œ��#�X��
K�)d7���KM�\�"���hb��ǝ'0Ź�D�K�'l?�<�������_??���ߊ98�=�Qt�yF87���@n�����u����w�'ޑpż�N��'��)abx(ʟ�L)כ�w�Wh�Z�S�'��e����	�5�y9^��Gz��=xn���ⴶUX]¥��kK��H�r����Q�?��n%,�\�WȻ3]`o[���nԭ���Hg�cy8�+�$��=�1�^�u.[��	vֲ���;�}�Y�,�������Y栫��Z� {�Mڻe��b��-��1٫� �&��B|���nk��/��?�],[�d[�}_��Zl���׼A4�n�<��v�:��H�.��k%��Ƙ�P5:xpx���\~�1Ю��������ũ�ڗ��'�~R�|i>�2B�?Ʉ@��ٙ�R�-���/:��E�H1��!�V�a��u���t줟�?���F�â!x19�/� �@+s�7 ��WG����9ΰ4��Mn��^�&��R�n^��a��v'���k%�eP�~�gf���8XT�E�8�,�C��׫T=|?2Tu�w��5)rĔɜ��g�̙�5��g���^��w>7J:w�R[li�Bu;�+�f�o�sm�R-2�  ��Øy�k�lZ������ϯ]M�dٸ�j�ڭ�=�[�`��y�鍔�w0M�⒧T@ͬ� ���[[��I�k���\�8@g�e-56�d��a�0D �9(�O���}�RP�5,��̭:��kLbێ�Kܮ��x)jb�B�dq)���h��LTeJ^�us�^+�(�i���Ew���Q�^(���'�jh�o)�"���8�I�޲��j"({�J�H�I���:�_�O�ss�x�����'o�ʃ:!>,J6�2HA�ŋJ��H�Z#V;�I ���3�t���܂�����s��W+�+ƾ,��PF�o�u�KdB�&ו??�i~���>{y��D
BWI�
]B���3IO��t�W��s��YCd�F�p�a�@+��C�N��Db���>�&b�}'�H��&�pT?�S�)���^2����C2!��Ǳ���!�2�!n��=/*�D<
�i����J�$�q����U���a���J.��.�@9�M��}V����k��h�(����p���m��6�K��J~��H�n!M���&�\P"ʦ7x-!�V�5�[�V`����z��@ �Yf�}ˋ�ϙY��B�4画@�Z���!��{���o�����ݫP�բ�M s�%�*��Փ{I=���k��#����Ẁ�&��e��)��cѨI~�i��%̑7��Z
ĤKǊ�+��=�P��i���dL8z��s�(2��><����p���� ���iD/��A։�e�D�u%�YiO��l�N�|Ke�p[@�Yq�C�5Ƒ<�,-�}i��EVn b��v�?rX�zEp�㘦��u�Sk�X�R=jW��IHS^{Zn��>d��.Ȩ��S�����l��ZH���u��T����Jf�#��Af�T�fO9����z�������_���x*5�����Cf��N�4�P���|����!t��l�@�3��+�Y-��U�c�����o	��#]���曏6�b�"��ݠ&����όl��\�C��e���1��}ݗo�T�����I
�`�;� J�gz��^�	�u^��L�YԿ���etǅ`s��w��I�Y	e쓁vsa�6�ղ����x���fg���B�P14܇�t��<v���b7!�D�-�p镽�����iL̀��9e���*��`�����A�KK�k���.
	��(7�x�֢MD���.~�ަU�'i��M��v�����[6短%���yRVsK1�YG߸}Pv%�.��O������_Ì���g=��-~���
�����抄	^�)�V8�Cz��/zX�5��J�� ��\ԛ~mK��6{@��6����Sdm>��I���:K��d�{`a0ġ�3 ԗ�V��hzG#�~c�B�S�3�gk��wq��K�7D��yU���][��LAQ��
��e��ಡ���H���b"ü�eبM�a�9�Pb�V8�.���Y��;������Ů��0�Ժ��H���wQh�����킯�H�%î�u�+B������:�U����N 0%�g�
I��,�����-8��b����V
��+Z�T���Z�[�OІ
`\���Z[�om�� .�Ki`���E�.��eI#�;�b%���z&�uwzY����/���Ǻ��yY��0�|�6�A���C�5R�T9W��LZ��oҿ:�ۈ�2C8Gc6$����t�)��݆6e��gOݕ�.?�v�|���3AȃHi��k��:o�F �!E����q�� 7�dRQP�fZ"&ή����ۡ��k�*'u�uQ�i������M5KsR���<�\��S�O�pJ3G"��y�����5�O�d��-�k�e		>��IGz�6�o�Y�W�3����b]���v5`����������@�Vz��ܦ��G��Ϻ=�|�sA�S�~3�gt�p�����kb��P��I$f�ة��������x��~�]C�\F��:���#�^u�70�\Lp�T��7H��a98�oJ�f؄:�U��I�*Ǫo���w�b�B�C!�C!\OtŐ1�oҿ0�A�����|a?���6P�`�������Ų# A�\�n
�ҍ|��7S�*�:�#�4<B-���71񦠥�������&�eUG�4c�c���d&C�{�X(�R�ҧδh/���� 7�N<�����Z��'�g����yO	mη��-�n�V|��~T����d���T�tť�"	ت:�h��H�nǊ�)ª����=4�?��@��o�W�fR7z��q��'%�欓V��9�z��2΍F������=�/�X�BUZW�O1�Ì��#`�����5��Be��xW����!.y�vvep�-ɏk�5Р,S��'X����(�YYx�M�D�5���e�z�#8t��tW�����k.��ɖ?bC�^)��Ӌ�Ȧ�9,�B@��M�d#&���Ѹ��s���m������=�_t�����@�G�f�#�����+���P~Ԓ�Qp�����
�Ϊ���&F�Vz�tk�����0�&@���o�F��ﵸ�N�	��y��f>�p0ұ�(Fs���lB�7fF�����7ӸW�ߥ�����V�\��HF�+��ԴOd�|�[��Ϸ�.#Y��F5m�]�r<�Wn���.������؞c`�3��tO+	oI��TD��` 7W����L4)HU�Ԭ�JPf֖�G��_����=���oR�,�q]fZSɱ�Sm/�TŮ��d|�=�T*��Jy|=<8�B�L��y,87N������Y�_�|Y�zh}v#6��J �t��s5�@�9�)���T�B�x�Ȭwv$6/�6M�H"Wx����:��|Ĉ��S���>h)|�w��ڎHs���"�}k�>[�[�k�/�쿜N6庵��%���W�g�aZF =�����!����h{/�)�$�͢]�$����0�9�۔��f�>˳�P��)c�7��`�IiJ���?۬���1���G��v�+��d;�#q���v��7Ybo�,��+��R��&1�|W@�7�5�-H/���:�$<�٫�v�A�Su���J/�yϢ���`��#���� /�I�C��]x��8�^+�ZY�i���*j(�eKG�h1����]
=|��z����C�^���K�q�A,�p8��`�8q��RW.���Z�ԭ��Q����Z�w�QYK�$�9J,Ξ��ª*���i�6,2��-Z�@J�i9���C��>[�#7 ���S4F��qED0�JQw��"�	iT���{��k2���"EK��e���BKGE�ШQºY����m;l	�x$��X!��R������3���ve	�P�e����������,8��6�GWw#˴��k�d��KV�����\��l�"�R��ܝ��	M CA�c��c�S��50�r��A�5��$�)w9&���W%�u�ڲִ߮Mיq�y3~Ee�@��j��̘<	_Hw�?dlq���ԩ/���[ʙ,�!p�f6�w\h(3�G�(���Z�n-�E�/y���q��_�'�#Q�O���z`]Ů�ꢃ�pH����eӅ�M����Ǉ��V �=(s��!�(��gt^�@s<�T��Fy gM��r_�w�b7Yں�+��G���̛�����[�x�;��~�%p�m,A!eX��ɻ"�r+��kr�n��:��硈�AC���K�S�N�QӤ]3l1�4J�[J������.��y/
�,��p1�! qk����s.�hN׏�7y�B|��܄c�Zޝ��d��A�p�w�~��+~�:.��y�j�e�}i�Y��坑��v�FT0�I��W#����Ư� ;B���K������i�ڈ-U��:�k���D��� GL�ه���@��MC����0�!�� �D����L��i����^��z��G�]cr�h�E�+'	���[�oi{���������\�~�-�(�JU[�YygK��r��_�q�6�&���hNH��N�[�-�N�dƃ2C��Ѿ�()"�u�$���������X�MWm��k!�C_{�$��#����Z�q��%��C�&O"E7K�#�֪ut�8!�IŴ���9R��H���tŕ�#!@浚��m����&�6��}N�v��xعdk˛?y��&��-p�X��6�u@�K��ϱY=���<!p��p�_O�i��}3�F��g�P�9eSDO�G8�qLh˓��x�R���d��jkRd
j6�K�$wA$��K���h��&��`�$���܂�U܌��Y�f�ӼJ��Y�#���I8@��%;���I�D"[*���1�c�ո�A�1�@���2Ԇ�b��$1[��6�Eғ�?�Ɏ@��ݿB���f�Ps�8� ��'���2M�݊��j�;���lCe���@�I|�S#
�!tC�h��Ӄ:�9�͢��xu���(�nڙ�i����w�>Pv_J[��Gz,9�r����֫��J)p��8���(8Aw��p��$�?�Kr�Ny/H� 鮷��"�i�@s<<.�ʏ�lmqk�c)�����Ay��m�ͤ��C~Zh&������BӬ`/�F+P����CiT�5�����,�u�$(�V������������۞w���|��T6����WWQ���5��\Ԅ����*Bx��Y�{O$�����|T�>i�˻9a�w���[^g��(�]��F�W���9��(Z1�;N�1t?>𨝽[�.�w ������TՄ�����j��c����P���lV�{|���W�J�Y�q��� !��z��@��]* x�e6�E��v"3��э�y���9&gk<�-�<���`)ӳB/Ge=�`�8*�%6ՠ�<�\v�������fL���Y��=5{%�w3�� �bD!���B�8G�z<⏆Я�E��]-�8#�F�*sH�pP�,H���Dj��ĵ�xo��x�WA�~7�R�y�4��["T~���6?Y�����-�*P��i[�F���Y�hk�B�P����[�*0�uq�U�]V��5P�0���`�~͊�Q��Xl��(�A#��|M��_c��W�0s�>{_=��" y���C�Ek��7�o�g��JE(���/	<�1H��=v+(2ɳg��<V�^�����i�L��Di/�}�������.z�T��o�1�pq��Y{��1;)5�����,��A`O �e1��b�\��OX���n8��I�L����q�	��n����48����8�N邋p�r�.�f���]O[�!<��G[vo��7�$ƺ��#�<i�2��z��2j�@R~}a���&eεx�z�8�.�W�D��֖UqqC��H�\�c!��Q�T� _�`𴤗)`>�}۞�4z�P�r{�!%�&�@�`¦
$鿵഼�ɆS�6k�Y����H��R������fa����P���ʀm�(
(*�h���Ή��g5�x�ý������Me��]d�y�n�xvg������=Z�R���c2R��E�U��@��ٔ���J�L�}��R��A�kA�I�X�#:�c0�W�6.�pݥ� 5ٗ��P���bI���j5E5Ѳm��טE���>=a-����vR�uU~�#��;Bt�pϧ
]���1���Cѿ�F�l�S����>.�f��P
�T
7��[�*襁c'W��t��]_�P�N���D9��a�p	GG8|6��tK]?ܨ2��K�\g=�q2���#_�bS��ɨxK��-՜p��%~t�6Zv8��Q�'�!��;b���/X��L\9nD�����׎&��ɻ�n|!i�q��b�������JC��U�Ε�!q6���e�y�e�ڨi)�(�7�[�n�Tq{�|�"���q���f��5��;@�Җ��M[�C�y_���s�ν��de$c���b�erXi�,��_n����i������s,M��N5�����M0
�W��=p������f�;f9^+��S�4� �'\���FM�Y�4pM�l��h��W�MN��-������v��Ś����.����,�Nt��Kb��7�G\�M{�dx��U��� ��}.��I��Ѳ�ʵ��U����!�F���������Yg~mn9X�=SY�	��|���((�����ʯ!���_N����E{˭/!	:�,MHxH����5u�2,T���;X�~�˧��o�X=sX��O*A\�{<�Ҕb�^�.C;�o� p�"�
��@"�)ˁ|��{R��u��|V���������eYQ�����1@�'��/�TM���U��+=ף�3���1�w�j����4Wf9���A0c~j�80'.N��g���=j>�=_� Z&RP�p�Bk�%���W®n����hbL���b��˗]�
(�q/�����),��	B_g� -��߲���0S�O}�!$P��8�l�dܠ�߯(FE�����%T1�D�����4��/=R��&��M��*U4*q��[/�-}Dn�b d<�8��n�OZ�FIBB����iah,����
V{]�ġPs�/����{uʴ;��RQ��gO���h̀ؿ��8��B��7����xN^r��	`U�5Е�w�4c/��i���Y�:396���o;�Z(=���r��P�p���+=�l+����w�ßV���j\g�
>�D�0/r��*mǈ�������r5�{����3�uǷ~E��ʸg �^����k���e�z*?�7��Y�&�U�kQ'���q[Z�]�9���j�[��9����^�m���%���+J�x���.e�A����vV�1-d�KE�G�˖T�6��m֍{�+(��S�~Z�2+j�3�?Rt�������h--J>Vu��ke�Վ#���$!/���vPCǜ)�yW��6(�G�m�(V��:�{�I�*cY��hy��(���g�6N��ۨ��������HP�p�`��|S�N��V O�^��d[�?W>^����xV������oc��9���GCiK�ן~G��rK{m�3���S�C�Z�y��yN&O�S��W�pA����?`^�_�Y����A?{���ڵ1�
_�2qӧT%TN���QIUR�J2?Ǭ�yC��Έ�iT"��W��,�rNz���GA���=���t��g;yx������q���8�����r�C՘*ks�=[�/��8��k2��kNL�my�WE%�Vs��>���xa��)5��!��4>R��L����{���Q�9,a� ż7�à;�y�}�+�G�\����0�\���V�h�ɨ9�]�<���Ħ�H	=g���f��j��x�8�+�[x���	Τre����	���/Ǒ�M���(�y,tT���K���?c'�&FO���~��a��~'Xb9��4n)^���.4�1�ޮ��i�������E)��Vz�v�$����DB��v����6�$8T��<��q�y�#��i�Na��0�Y�~#�m8꘶#R�~��GW[G֞�iǜ�yez�0}�%���>���<*�8�3p�uXk����l1���p��s�
��{���t�G��I�=_£�G� ��Ԅ��H�j��np�A�V���]� O�V�NU�[�}wT�#X���UaT=?�-�>p��g�ZI��"Y��q��Q|�~nuJ5v�|��b��w����E!�&3��`E�W12�?>�c	({���Ƴ���M�܀Ǵ5�~|��E��Y�rD���ѰTr�%v�A*g�7b�w�J��`������O�v/�z�����b
�c!����A�h�|x�6�}�x���X�FJ���z}�i�80'���}�D��xq����VT��~�G�� �e��"me3|0�W#G���^�� U�-���D�����y��:D�v;%�	1pWY����6E�%#6q�@�?&��V���]��+d���׭[��$\���`�m�ON)A�0�pwK, �p�8�Z�@��8�j)�T���-�1���L�	��"p�ޛ��{�~K�2����=/���/���Hv��v����BL��o�P=N��~�x�%�U���h�����W8re�(�N2�C��S]�K(��və?��]]ŵ�~��
��iWK�Z�U2��ROWU پ���-qR��{��޴�dw�:9Q�|[�x�֖�oO����/`I����Od��&��[��E�)�x�ȍs�5�nU.ZoT�A�j^��|>��~ f�i˷t�ZJ6��֮��4���?ĔK���l`���HS��]�Ix-������}�*��-7��ج���5��i	�OK|e�z!�zly_ߓ��n�&p���V�v�Ϡ����l����cPmNw��`�v�e(���h&�N�����W[],��o�4�bfc�f޴&��Z>�_i�;��Il��A�^!��^|P��i@)S�r�F��"&g��O7aR�<�8��}�W,����H^u)��?6�=��X�쓌�/G�[�7��]������%8�ٲ�M���)!r��o��臲O"�N�%O/vv)է�X��5}����g���h��d�ب/��v5��6��TmPk0En�o�o��1[���8�<����"5``R靯�$�3ql=������_G��S2�R��ۇ(Fp�rm�NQ�>U} 1�0�����L|*�[��ф�ڙ:�j�v��k�=q��$ܵ��p&M=���*AvBZ���>���5<7܂�Z�i%P��4,�{�99>���S�7�y�X��+���(�]��F���^��p���]БF~uy}����8�y�+Ԩ��+�B�l�)�"���3�� u* �Y����2�S]�_�x6���4���ژ:��L1њyineK\�ھ��̻Q��	�����]��?�tɬY�#N_�_F�s9�ŕ���;V09�?�2N��;n�	;�FQ�҉	�9��d�o_�<a�l���ז
ٽ�]�T���B��D�4�M��QNF�"���G�E��" �	e2c6�?���/�u�B�.J��'0�W�+���s�&�3�$Z�"M���� ݭ��h����X�:�8�w���K2I˃��9�̲�6�.S�9N"�y��<%;[oqSm$�t���@`�={����X�}��>�,�d/���Ã���W���n��L%PT?�j�nDK�ํP�y��kQn*;U
ㄫ@�2BN����8��쁾
2fZ�#J���)Vq8&��3W}�*����9r�˕�=1��64נ�6�E����[[w�����8?Af�'¦��@qW{ɝB
h��r��� gGu�}���U��AL����!z���%Q4��;vw(�iy1�d~��Gm�2s��ĕp��IY�dڕ����vAL]N`�|����8G�ao�X@}f�M}�~�Z���X�:����`sJ���Q��>A�n�	71�D���ر��E�R8�\VSA?�Y���촇��E�k�G�3�|+�B��$xn���|ԛ+;S]�/+�@�ȄK:�X�_����TV��T�;TL(.�#��d�=�q^�g��i�����T�x� ��. �#���\0���%�� ����Bs��/2����,��̍NZP|��(nD}(���+�gg�,��B�6KN�Vg܊�e�hJ�C7��]��WՔ!.Y���Y&t��`mrpF&{F��_[x�f���9��)m����[G���b��ntQ/9�4'�hW��6������	�D����X�h���y#��\$Za4?g�ߜgٕtߢ��_�K�b�B>�(Ә)ĥ�|,k��ҷ�D>N^�V=ݥ�[t\�Aq���UK��çp��x��V���w�'wŦ��9�q����!�i|��2��t��b�T܋�U�9�9�C�uL;��3y*e�Z)��ɼ%��}dٲ��N_%�	��E ��n�Ӂƫ�C��d��B��U{�y�آ~1�{19<�%���=j���k��vu5�m�$�f���E{�	a*+`�͎�q����U�Qh�)����(�G�m���,"�/�2���l��[��FV$!RJ���0���'N�b= �n�:E��a���UpSKTl��"7���!*E�!�������)����������ַ�5��'�?�¦���+�@�D�3r�\�U�`�M��7{��#K�g��q4� �8�al�v+��/����A}=���	s�=�,�o�ѯ������W����Q%�Oq��6B���nR����Ir*Yu��Sn����Ki'�����Y�K�լw��Ŵ�lrz�.���΁n]�j����I�9z�M��P_*:�=����h~����#����J~L\��Ph�ղ����%N�x���E�fJ�\��¸��� ���r zS�j}f�CN/_�\Q�$Fu�:��h��՜%^�y3ĩL�j�7t�ϫ������l�(q�%���S��Am���\��
CtG����M�8��b�`�W��CB��h�s�̑�V��+����0
�}��u����ۡ�CټX͜x�,� S"�6�*��6�{���7I3n�� ����>Xq�k��t9���*TB���g�1U�}�k�����s3+��_Y�e�_�=)0�hi#N�gn�]���a�<bj�l9Y�"O`ڗP�tH���E������=��7%_�fOG��� _�gH����I`:gAK���
ot�Tګ�x�$�n/�gGt��,��HД3,�-[��]1��$GF���*�A�v�%�ќ��Y���p�)�Uī�">�O�R�n{O�!21؟a#��D��pM̫]���.ya'��)�m̘|>r^�v���"n�x!�ǯ�u}l3I[��Ӥٲ���S/n��lN� r�0j�k�R�X�U���y��q���DJ�?^����C��4
�wW�Z�\�"�:D�/g�#�^g��īv��^csx���CZ��Z�PқZ5�@J���_Km?f��Ř�Yҡ~1��/k?�DS�(�
�b�6��y��U�%�n�J��O�V6�����J3��ʄ���N����F��������?��X=@�<�i��1*Y|PDS�N� 5~�k��I�����loli�6��xv���*2�7�?�p��3�o�<;F�S�q��z*k���lE[�G��E�-���ZN�N�z��:�~,�|l�Z#�O�G�C�>�C�}`m��+��K� ���#�L�yPťɅ_��C���i'��^9
]3�3bFG{�>��=��\�K��R�M������rr�,�(�f�M���HGl����� |0�\�>cZ>ͼ�`�2)�αw�͕���I���_2<c>_�I���64[�g���&�"��i`�$$e�n�2�m�L��t��� ��$��_�H7�j���; �#��JYS�|!_�ql�~v�=�]�3�S@4�s�7������TKA��=��a0w��H��%J��hC	�~nF��7��u�	�0Z���ĥ�x����0T�����͒�a|Q'�O9��7[	p���͛]d��Iu#�O%ˣ�L�����aM����~P����~���0��bg��M��fg]�?w윕!����X��љHi�Y곐K+�k��9�IU��hm�Q� ��J��L:�$��燚�I�@u�����N���*�|�r^�.������[]MZ�#a�X�nx
��=�!��a�u���
'�qA۩x��>zvκ˗��@��P4xÜvN���i��'��K�S�|�K%3^��̗�mb3����a��ʰ��M��]�)
�KgԞ����T� �a��ӆ�q�ҟֻ},��'b��-,�����Eg���B0�� �%��e?&1�6OeA�8����p���W ����h�T�36<��F�t��q��W`�a���E����	���Q���B�:A��<���S�
�kG,�{}��ӫ{��?_ �j�HzQ��*c9�+���5Odژ�r[g$����^׎�l*N�P��@�$PY���e͆E���"��J��@*Psc	�K�`*q=I��\3,$��<��D�������X��4)�A�E�Dp�R���|��f��^�&������X��CQ��\9�,��fY ӾK����rp��4�V��zP���<�?���ZKԓ+�Y�nDd�St����� ��)GQ����1{�e��>�"Dz�}�$�!���@Nٝ0q���!�7�-�Rf^}2�r"@K�;�=�r�� Ő�5�W��Q2"����n=�ydBD����0`���ڎ��$�r�Aq�Qԣ
�uw7��`k}�!.om�����4�?1��T����:y�\6���2��F��C.��؀���և�C㟾/���V�a����nyqgF���2��#����rB���<Xw��"�C@��Os�䷗���A�#ξ##������m`����v@�60�`t�أ兰�21V˦���E�̯<&�9��S�+=w$o�R�2�*!����L2K5���GX����O�7x����R�I�Έ�-�~����$���%�2�g��K�6�y��8]�=8��r����ƒ��E>Au	�4��,�XYiB4�k����-���a�9���Z.�G�� ��mCR�Q`���d�?#�n
�O�/֭$c���R���-[؇���M2.�RDUDq�n�ْ ~�U�ߵR�fb\�H�Dv�V��PJ�>��8K��{8��mGKD���C�1zk�2]�U�[���uE�w���G�@/Վ��]�	����Av�f�c�.o����F�˕�d�9a������r	�|���{���[�,`>�K�EE�**� s /�9_fD`E�io'�����/���
�W����_V�&�� ��
�ǅ�B�*���_K��U�$���g�?�����?\�s�9]�#��fP�+�6d�OȮ�������UyQ4�{>�V��R,��SoR��>�Y���)ΰ�!���~���֤4%�@�#o�ai?Lr1�r� ]��&����Mu����W�ĢMVj�g�>:L'S-��]�-����aҡg(���gF����K)���&7�k��ϗ�)V���.�c�G!t��E2�	J�ҕ⟛��'�7���uc;�?~�\s�8SX��M�WA޹]����g!`V+K}ܳ:��47tX��O�f=��0Ԗ�X�q�$�(@ʇ�R�`P�������ڻ@��@��>�I����߷��ol���n��V����$L1�'L�~tMry:����+���E
˄

�V
�
��؈�q�L�=�r�iB��N�L
��^%U�#�՝��,��3�II�
{��5����VB!Ov�l7�Q˚~� U�oL#E�
���G�H_��ʢ�ƋJ���kA�#u�{Aj�F�'��n����o���Z-�'`T�[x��ʴ.������A��4~���Ӓ��~�Y�+m�MߵD�՛�fK�ͬ��5���B8��@1��5��1��~Lz���S��+nwȦ��Ҳ�ٌ��f<��D 0�j�Y���>��ZF�1\ޙ���Ѯ,Z�^�Af`��]�ȥ��@&j�ߕڀ��:wf2ζ�Ei���Q�(QO0$`��� �Qm{0!^G�0�����'m��|]w
�_S�����2���_�U!"��`<ģ�
Kt��;@��i�?Vu	�k��&���Å�/5��oE'{B�[�i�8V�8>�i���W�`N7�N��i�a��)�%^ENW!�C���u\�XD҅������gm�X�̟�v�d�G��V{ƀK2��C#��@���Y�'�I�����Nuvʈ~p�iz�!�$����weF�V�jk�;sT��,��j�)�k9�lBo9`��Sw����|�� ��+��W(�p��+�ku~"�H%�#t)������[D����@gT�ӘN�$	N\�M�϶M�a��/������(K�G�Q^L�?����y�]#w��k{�S��d-���!^̬�&s����Ǉ{�D�F�%:��g�Iˌ5�����oI�|}��5�q�����L)<��V�q[4Ѕ��y�}�ÇaS�����c�8��#L�g_�qŖ��l-1=�
b�H�oܺ��K�}0�&�M��V�F��'~��@U���oR@�De���ތ��{��o�̮޲<.iG��G%�	��r%����h麖�t��ٓp<��uWaz��X��u�e]D����sA����%#%�o�1��������`~��YƄ�lգO 媤�3U��ywg_[�Z��4:��)x4T�5����$��Y��~���r�K:��i��ֽ^ %�3��H$�V�a��(:綆˾��l�����8z$j���+W6�rM�	�Em"<t���A_}�s��W&�O����n��d���!	�����.p�A��B��}qD�媅,��ɝ-fK(JpI�e +����<�"�f�ҝ݀�����Kj����t7:�v���8U��]�:�.Fh^���y��ɟ�0G�s[�aߗ��G���t�䫶�-��<�I��.�d�}��b��_:F�Z��&Xj������Ń�W�<��+cGG��ӧ1fM<��T��w[��Z�h#�ļ�O.�>��\V?8R���=.�n4E@�ڃ�]aL��
�_����������j��Vk�7F x8��P#h<�·C�K����E�w�Ae1͆%\�]i���P�̻��X���?��.�>��Q�� <,}�˦��Сk���<,�)���HJ�E�L 	7��>	��?����P����v�P��	��%)3=��+�W�x���Q3>���"��¸�f2�i��l
a�fp>3�����.�sK(h���?H]���e��D����c��%��В<w霥�fGlƹ��E��UE�!��{�GT�P)g��
ӳ��H�X��O�aYT��y:�d��4��JUeE'������ť�� ���d�V�>ְ��N�[��g��xkj�W�����S���FX9�5�l؋\��4%�fi F:�p���
E*���rj�h�}2��Ƶ��7�nT��ԡ0������k�ܾm��P�C��%)[�����=��|� ����@$G&kk��6��!��~��!�!���%�����N#����z���{�8�h2�cD+��t[�vG�Ps@Ng:^�6�!����#l��%���*F�8[qn;�v����i&t+h}�4��腫n��}�eߦ"h� ����ʲ~&'¶�5 ��{��$~	�RKvc��C��Bځ�a:gG�a�5
���О���3��uY�y8D|M�Y�����7Ȣ��`�c��.��7��Rymt��[ͭA�*�J�r�@x]��jB Ka5��Wݞ-L�4.É8jt��0�,&�F�Q��@���dW>�ƺ�3L�X��;�O��L��wV��E����y��1Y@��s��.��,0�r����,���������t��هzլ:�mƅ���x�ZEZ�l��UV��%]JL��Q9��<�E��1�y��&'�v#̂��2fƞ��i�-t��N�6��:%N=ت-lG?��?H�>�k�<"0�#i�����8����7¹~��.�L���
*�UTш5��CJV��)��(}���h&!?2�~���/=��yS#`4���C���8�@�/� �V�	�B؎�1���6v����-��"	��x��M7�,0amt�	�psx����w���'��6[�1�T�ۄ&��;���1�s7��L��w���*�RW��-8eF(9s�.�_2��.b(��ͪ�P���u�ah]�X��>��x/�m��{��?,�I��E�Dm�|˳{�嫒,�i�3e�O��y Ot��,��V�������2Ylk͟@�/(/}�4W��Q�)�����3hC� - �1|]��� ��sp���۠b��c�jǉw ����`���N��K���"��s�44��Ԇ��I�ê��J<],Q4��>xt����#���Q�5�H ��O��pJ�ܷ��k���h@�#?��,'�V^ ���ɋam,�_	S���Z�*te�wP�L����|�\�p�/Y��a���#%��.�Bz:�((��?���H��Ķ�gf�W/!�����Q9p�k���#����f)[r����l�d�*�C�7�0�����t�Cz�,��B�̑F�8�7�=n����;ķ��g~,��7��Զ�m�$����%㝹�����Z�����Ό�#�|�fA9�1�щ�p����lDz�̃�)G ��ݣ��?��xW�K���;�»� `��b�v쑴�<^��i�L0����u�ú��Fu�7�2�w�Z�y�7�%���7 ��=2<h�rY��3���4�)B��"�&:��h�8�e���m<������c%*w�	F�	1��i����� ��ߧxυ�up����ERt���C�dq��,a�$��#��!4� +Y�iꔽ�;�HF�ȳ��������R�� �Q��[M R��=N��R_G��w.���Kʾ�荇8����&�5�8_��C���&�NvSK`���Ǉ��,CUiL���W�g�%�8����ä�,�9a���r���B����Λ8'��3M
�Ŧ�1z%*p���@��LnY�Ϣ�e�z��S��l;�ѯ��-���7�nfDN��:7�'��5���/�r�Y�1l%��cN~Em�w,���WU1��_����	�]���oR���j1�:��6"	)6쀏��5�c���>Z��q$!�+#��d���ya{˪��!�xx6F� �#M���l�cmMzC�t"�k�[�;^n�>��8<�{	}����60��;�L;��{&f�
��S�l:���c��tz3����jy��@�EA����G��W�/��k��ݶę���@G�e;��6�3#_�)���!Uř�Xop%G8��EZ��"� �;�5N2���
-TtQ��ݘn��1/ct/3��K?�����` {M����_�:z����VhH�T�2�eԽ�@铍qg�c����$�]��yw�Sū;[��߮��ft̬��N��H�to{1�\�@��� �B�,�Z$I%{��/u�&��iB�*�1����^��Sc���j���";��=`��\f9LHo��ܑ ��st�I�АR��x��ͧ߻��q�I/f��&�����P�W�V�$���it�
ˍ�� |��%M�o�Fj�bJV #M�BB��TC%,�;��:5�b���eb3�� �;-0��v%G�RK���� YZ�,�$�C��>�A��X�m�(�_�����F;�����γ2)�4���zI�6M��w����M�:ϑ=<P�IK"-��$��#�(p}1�l\�n?p5��*�?�Q�8�}����� ���zm
�s!�F��~����P�5pD@���
�"[}j��Į�`�����h7�}j$2��q��c��%��d���B����[���Őd�5K�������������������HW;�g��C1'p��ݤ�Z1mre_����W�1�!w��������D�e�b���Yƃ��T�"��������b�4�K��q
IP��U�� �~ȑ�����K�Ia���cK�L�*�bLU�XR�].����Υ�@�����O3��{ӧ�N��p^��� G`�*V�H��\�jqT�4+߷K9�j$���'D�.V#r��`�ur$�3�0�S֝��b���{j��r����d���^cM�nt��kx��'�6��u�Q�G�V<�����]�ط�(�2\f�[j�ǯ��f\��즣�p�8���ϓ�'w��@�D�M�U���j���]Xb�J��W���m��@��	��3V�5�%�,�#K&��z��^u� ]uioAȐ��7U�L_����25���O��GPu�h�����J��������XC�E�����	�.y���Gv��7��-�0�5"Vo�c�^��%^ZaO�Ŋ�~r�|?4�����u]����s����޼�gTXS����B�����y���`0u��(��|��	���y�$j��������7�W�,�.Q��!��J��QE��]iT籔2�_�|tR.�B����d�� T-�`;T�݃��&Z�kG9Aց����n�c.M���H	�Q����4[�D�7��`�z���RjD�x��*�,g����~SӮb%���f.�*q�^:��a��C1!`��$(�/�a9���ݼeWsꯊ�L�.-���Y��I�ʢȽ"
�|� 5�!�1�B�Sz2������ٲnUgD�^��krh��G�M�
���ϳ-�zj ��J]�$��'_��!��盩:�g�L��>/��Ġ���\*��z�Fv��u�@}����S�;�F�el��/��ڼ}Rh�o�P�Q�7���L�<#��4��.nSH���y;�5�ؚeډ��߅c\�}�0���cJ�v�Y�]TX4x�����.���w�yQ���C����o��5uC�;F��y��Gbn��Ʌ���ʰ�:w�ױ���(Ϟ�]\������\�Ʋbt����	�A���B�)�0��wo3�����QP�dې�_���-����~�2R�%��K
�����#IS���$'�P�U�uǉX-��Za�]?y*��^h"z��.�M�,%5�7���Xh~��Tm�r!�	.�G��&��D}�ǜ UNk�U��V��&o�6�3��45�/���=�0fu��&J?Z�2z���9j��I�6��Yw�r�(�^�Co�g��(
�,�tnhr�s+��;���{��^��MO�H}�#�z
N؋�g0ͼG��~���K%,g3��M����^ǿ%}�X����qu�/V�#�I��؃�uGq+��e�*��������g1��U8��-���IZ�?��nN^�<���0ɀ��Th�JoϲO�'�`��ơ=�П��Lt�LC��'��}��|�D5*P�ʇ�Vݤ�z\���.���,8b��@B��o^I�[])j�t���ĵ�!�����bJ|!���O������٧d�wj��%%q#OX�U���S��^�>�IM�Y6ь3������r�A���y`�XC��V�}�nk�h�e��l����Խ+�"J�C!�n�_7�:���3mH#�%T*9���ǢxW�=�l��{��s�nS���x���&��P�i�rw������߿4���`~w,�i����MOG����ys�%ʴh�{3 Қ�Բ|"���e[TltO�g��,��p��ZD�<9M�O�H���!�A���Va�ub��ɏ�3�Ih�W�PE���(*�GR�
���\3��cq���n�G�
(jf�����ϻ���7Ɖ<�5 ��F�IЉ��X�#��r�Ϟ�����w8P� 3��U^��z�͓rў�a�l������'���ֿ�d��| ���nP��M�'P����F��������������3�s�-����iC@yd�"�F��g��L�%M>����)Iz=�@!9v4�B�r�_�[����nz� ���̑�5=����cbVRmU�&`�
�q��`����'�K΄�)�z�٥�7��G�J>�LzV�3���G���LH��r)a���D��CV�e^���=y��ż�ෛ�2�C��,&q����R��!Ԫ�΁�b�B�q�I��_3璿�l�؟\Kyq�+�nlo;��(]%3w���.p[�d7r��)�´a��O/|��t�C��:q�9���X��o�,Ҕ.���N��ONU,R��1�Cl���d؋�����P����t���J<]-�J��o�y����ϲ�h�%�&�ջ��YG�KD��H ��۠������%P�:�B�C={�� �2��[.S6o�RƜ��sN~m;7�Q���ۏ��Z�so�@߻'N&̮�G5+G�u:�m6��P�����Gu/�/�٥n4Y͉-�}Y�
���c(����|!���!���@d�q�%י$7�����Tg>Fvж��3����z�����>�~���B@،�!�Ɗ�q�z%H��q��f�&j�pn]3ȳ](# h&��+�,�em�/���&�=-�r�[��G�יm��#�����Ȏ^v�n��e]QQA��"�	ԯ����W����!�B�BW}��k����zKɀ������_ID��{7LY�ӱ��l��s��p
�c� ��a�ï4��.cv5M��m��5����4�G����(�6-��R����Bzl7�&$GR���:���Ǭ����F��t�@uC1���y$���d�Кy������8��0��c�ҕ��`����0}׿:�<fY�_�9ޕh��z��Lrp�ןIG��9ګ��
��N��-@yH,I���T��ܾӇڼWL
?����k����ƾ+�0FE�͕3)�:�l�tѨ����y֔�؟�*cŌR@ŲAܡ�]x�bf��H*�4#��A�Mm�2]������Z\��)��-{	)س���lxp'�[Q��Ohv5k�<Y>U��e�w`�0���/%B�l�'�e���)e�Il"�s��QBS�����-.������_sgLd"&�6�5v���m�@�n�#������ʇ��ҷ|��#Ǹ���������Hz ��B��T̩�b��O���s��h������6Ƶ9��
��f�ڦ�@v_�}S�b�0�q���
�*Ԃ�`��l�Z4����2�5��h��r�p�w�|z�:���yM�:�7�y��E!�N.�At@�Dȿ�b�l��O��覀"�ŏ�"gFH�N��P�2"s��(�z�q��=E��}�t)$�H���s�G�o�����Nǋ��2&�����-�fY�<f�	�nںTtͷ@����6'�.�a#K�v6xqR���#���^�q�TT�9v�f�0t��e��c��x�:� �Q�2�����R6N�p����	��u�5;r/�B���@2���_�2�Up3��Q����*��S���c�#E>뜜��i���:u��f_'_�$�
dU�O��4�\������&JN��'= �X���I
���jR�l�'SK`u5t�jJ�'�`p�u����d��gȞ�sd>�t�M��Ϗ�	Z���[[6�7�f�r�R#��;h���~M�|�>����K�U9TB�g�y2X^�U��/2�!��1�n3�����DQU������
)S����4�X{��j�cU%	[�b��v�گJ$�i�эN����tO���@�y'bz!#T�tWra̓��Bus�X�>��u��p�G�U'g��q}��_��-N����-�'� �K�x�
q���a/*�u3��)�-�5���њ~}�Ѿ-(�4��˖
������bNi�Y}�k&�M�'`d!D!$��}\���&5�>�:�H���yy�f��Y�T�D�}u���UF!�
I�?;#_!�=$�JD�`:K��X�ԦQ����Q��ݕ�C�m�4�MV��-�p)�{i�۹2t��ItZ���3q87�����̌;3s�C1 �V��j��o.��-F���|�r`G5���V����iȞ�z�֍ZR�Iw�?"Nm�{t����,Y\C!����:��#�\FRq�\}ͷs�X���/���9�#��[e�\�hx)���?���F%W�:W�b���ٙ�� ���M՗7Q���G�d����6��D�E	Fq�S�~�j�/��Sƕ*��̤�\`j�G�w��2�hX��`�����
"}���I��B��	J���츶�|�����3ސ 7[��b�_��҉���ai����AC�Nfd���e�?���g'G����@�HZef��8��,-a�S�jX��d�Q���iK���g�z�'cJ�^g}�:�.�`�:^j[�x�KA��G����h x��`��Wn�8եu��0az�+�جG�#��;�����wD���i�t{T|(:\�49a�sKou��P&�.���}�9P��f;1{�[s�Ϡa&\;��]�y}=Z��� /Υ��y��js�辿]�OK�5D}a�����9���XG{8AqF{�k6�ǓՉ�mj&چ�O*��B2۴�Aϩ�9=f�bO��t��RM��7�:��ſ����C(�7--��#5���G؄��g��P��|˙q�Y��q7o���v^��������R��ND����/)"�R��3s���2����.��ƛ;����#_]��[<򗉪��v���fҞ�P8������g<����/�=7~z�����_X�8��[�O
,\J(3�:�n(o��*�m���6��]K�f�و)�����d3V{��	��RJ�����α�M�޽-��Y��OY�X�s�1no��t��^���8z�4��Y5�=��y�OP�T���v�����P�ɚ=ꞓ�-N��+V���Z* ,�N�x ~Ek��(�дG�S��Uϱ[Y�>�Qu�,�b�t���G6���!y� H�u��H�M��w���8-�>��oT#���J������ͨ&ɒ#r`ϣ�����UE��o4��6��l?�L)z�5}Y1Tυ3��?,��˓a��i��W�X�{URD���k�|y�?�&���p��nevF1kc�&g�p ������óV�/���N��
�ҌC�*2�w@�����cr����]3�5�0�>�2?OL�4]E!�G,�rJP��N�=4YCO*&�6����P��y%r�/H���վ�W�)ʳ��g��ȳF�oSl�P `�����z1�H	�!�rF���dOE�/9J+��-�v�ϰܕW��'!��C�<�O ��+)�ҿX=T���%�T6�v�ν�?��7�"���÷�s[X���4��
�_��:0)��z�4D�R։���ښ6�^�h���)�c����|�FsEosd@�
��hBd]{��M��4�}nnhNVy�ľ�C�ϥ'�G��h��$J#i�]l��_/UөQV˟�6��ڔ�o�Rj��:��1)�z�`�?�^�l���!s��SB����"�.q��t���ȋ)�*�[��|��cL*�G���^��w��T+@��$��
}��Dfִ�.
�w�V3���j��;� �Ԙ�Q{��]I����hx�^v}��I%�X,�CV-m�I<�rl��D����5կ���`�����!�tG�u]��{7yt��K(�S����[���0o!�I��6�����&�*�X)�Qf�$j_�qq�݋1�T!1��q?���P�<�^gu7D�c!5�o�>�iv.�hN�fё�Så}��|n��Q����G��� i\��@W�A׊�	:=e۬�j���Xy���K��R!�$XgL���V���쟔ό[�P��r6yT� +(�����S�%�M�岐}����*+'U"p��m����,��q�"��<����ȕ�t�܊ᔝ������ذm<TĂ�6߀*b�-T(�+2)�q��5�U��dݭ&wƀ��O������\�G�#�����~�K�?W����P�*���&i�U�W�b��,����E�jV�ސ�	)���3�l��rwÄ���`TL�t�E�Z3�{sw����r��m�	@덑\e႗����oʈQ��i�d6UJ�l�Lm��}����x�2�kM�ȣ/��B��@�H��EӨI�m��0���o������Ē˰�R��M0]P/��+��c���>�LSy�9�,�4�+v%��R�������l��y���e�>}!����hՉ��%nh��R�b��䄡9�����>eI�|���,�s��1>p��@"�bۃ�r�<ml	�9��]�#�KOө.O�<DM����U�;�K"L)I(JV������}]-D"��p_���jp!ľ��������Yg-���%Db�>&��_�<��ɳ�k�.����q5-�-{�_Y9 *�/���D��:/P�1�Be�x�������"2C_ߏ����o�� �j~������?�#��M�S ���m��5Q������?���E-��+!�*�t�R��b��6��LQP(�1m�����|Ӷ�5�-6�G(c~|RB���X�QL���P��W�W��!���䗘��6����p�ҫ�]��2S��C�r�������Z/SN�$���`Gteh�T����8uw|8p�Z���]o�c$=���T���/�և�&��ܖ��|GZi�A���k�F��ϱ���>��6cdF�������)�7Zߚ�\�_�����K4	?�=�H �[^�7�J�.Pt<�Q$����'�3�E���2��i�|8@��$(��LS�KP�R��Բ��g4Z�Y��!�B�)�H)�j�c�3W�N4�.ɴ�;���)(��8V?�q����kw��x
,��ǧ���֑R*���^��}�_*��������A!��)��d��9����,�{8��a|�x]Oɴj� �J_B��x�Q�l�#�*��&�ia��_C=���}@f���`i�9knTȍa��x��aZV�%߹hQ��|	K���	�7N�R��>�C��#�c>-gPӖ���Γ�U����o�@�j����P߁�`)�:���g1����}�,6Β��P�G���ɦjR��Tf64F��N��B99��YB�:f(��
��ރ㕾eTVfwX�jr<�R�,]�]+\ʗ�+���0���?���|ɲ����䶈�`zd��Ƀ^U/"I��Кl��$�Z�O][^�"��b�d���"� �JD;�dhٿ��Fd�fdTv/��ѭ%Ca2[����K�J{|Z��JOB��7��X��!s��*�-��ף>ۉ\���� I��%Y,��3.*餕pd�a��ڻz4�`Ug��{|P���Cq��\�C�0��Q��)/Z�q7��ˇ�4¢��I|-������]��A��w�"G�����:Lޙ�H#�-��^٨eE�� �uG'&�]s&GIXɶ.'�0-�&�w�r"�@&��(�f.�\��Gt�I�X��5�����ao�d�s�{�r��h�(�D�7��Jv1c�<��FE��v$��g�@���/�#���~1Wg�2g*�ji��ʱ@��*�1��Pyh�����O3VO5��E���w"'n`/ذWC�[NeF�k�r�O�>QͶ4z�A!�+r�������dh)�^u�G38ru��3h�m��6��j��F����̥_�/h'�vy5J�x�.4� =���@��AdbZ��1�0�JM��0;�u��Σ*6��~�C�x������',g>6#�c���S��D�[7�RY�?9�ڸXe��Z�==�p���C�v�}�{����Mj�r�h�bj�\'�pDޯD:�p7Ѕ�=.��yK8����A�lB�{�n"+[�x��`
�YT��BT�h5�c-#+��c�?B��
�F��-c��|�_���V�WF!�|DL2��ׁ�a\��{{��5����>�z�}��)���-mi<�<�땂(���ry��x�p�j�廌$�ӧMM#q	�s�PPfIF<;�@v&:�m����n�
��AT�Zp���`��H�ل�1�s���ʗ�G�vR�Ɉ���6��s2J~T��d����{�h&�G_���#�72��?5���<��!aS�N`�wu����l��ҏ'�;T��QZl�7�J�Q�5A��J=���i�Юr�mԇ6�ŕc�֒��Vӣ����@K��e8���4;-wk!:t2\�����cd'r��~��S��2��%��]���lk 8��!�����VrA�e}##ߪ�}�"���(l��C��M~��YN��'�r�!�N*S\�Y�y�^�س
�EN�h�m��/����率�y�x��u���ΜS��O�9����{	k���虧I#��\N�rFedсx-'Yj��4�'X\�Opn=$ro+Ə�0_�?,���P�z���0YJ��� 9D[�����/��KB-8d}���L[��#A8(�̀ۉ�<����)��{�$(a��k;�z'6���4T�1�1�'�F�����{��o�8����o���K i0m�fN��]j}]�?!w@v'�B?�6ޔ vkOs܉?�~�&�+i\ĭ���M/ꏹ��2��jaJj������`cq���T�6�v��P�/A���x�B�.�gt#x@^�ȾVI�!�$˧P��?6�huݸ(�p��s�Ht�l$�����)��O?kԘdU�E9��'�
�5o��&�ŝ)����ĉ�2	�À��4�����l #�M��a?^��I�Q���&&rL׊���Bc�]'�G`hZ����h&�툂�8�������!w���]�e�y���!6���]᎕M��߯8�,L��<^L��G�n�KPabG��1�hT�5�Yi��4�i�o�5�A'�,6��[;�Y	�I��,��b$�`��R��6��.��z[5��>\��s��i��!]���PBԇl��s��<�:�,VT�fO,��8,W��C�������J�\m�bv����6ı
����r\�	�v���\pEw*H���;���vJ�7���p����^�9�4��ʤ�I�!�M-*7��t�$$d�G���N +jz�VX�=*�ʐV��M�Zh��t�|*�?:�������N��������T�5�v�
��Ջ�.S��d*[\�*d�Kⶼ�-��ч}�0����>�NaP6ˢ�� ��%�ș�a�ޫޑ�3�U[@b�D���7~\8Y��a������<�6ᇑ:Ǖ�89���W'J���.W'l��d��nG##�X=�z$�d-�YƟ��!�v�˞�& ���WK�)k!z+Ѻ��4{�'i�1M�J����I ��g��w��^�A�[H��
<.a�+����b�Bt����7�m���B���R;�p@=�^]c���)��5~r���SZ@�� (�	��!�f�^�0�be\��hR-�S�mg��=�C�2
\�p��K�Pq�K�p~�Х�Ϟ*^&OO�i��G�Ib�^�Q��V���e�?�&/�����W�C�^�di�4�u2�m�3��nOZT4�\{r|�h7uȯT<�\dF/�b�h7N}�ط���l�L=8X�S(p��J��bl��ebڊ��m��{�xݷp>8L��?�S����@���H�JLB�2�x�<���h���[���`�������X�B*v��ԁZ�_��F��Eѕ5+��9KM��9V.��z
j.I�Nf��TYL�!g/�I�
�%L�>{��Ӈi�}{l��ia��>:����P�.�E���]a���m�-�I������q�ò]�Vfv%lT���s�i��IB��=V��W}x�S�}�� �u��Fl|�:���D�����̷C9Չ�*ǀ�Ne��)�T�[�`�խ�Z��S��"6�}���L��e2m�W�������%�
6��� Z�@z�L'Z��AՒ��r�(���������}`Ҁl�N5{t<� -�����A�O�p[uT��@�0+d��R
>U�]�4pD|~�+ja�����N��y��ͧ4 �#ѹh�H��+�]�O	�C�3����V�d>�s�$��>~����>tpǂ̗R��?�p�����D�,ᑫg����/�+ɘ�[	4��-��!��/\q�(��yt�}X.�����ۚK�ݔD���H֯HkX�x�]U�6�0�^�3�!y������Pݘ�ڬ8��
=>�Y�� }��T�(�.,�W��M�}tt38�Ǿ^I6�b���4R1����K���Lq`���ڎ�!�Nķ{��)�X�K��
;�[FJrK�p�DV^��3��z��������2-3M��۫��T�YQ��]/Ŕd�	���c���^04_X�3�]s�'�� �7�a���e��hǊi�?�.>��	q�x�B�%�P��.҂cX��,Ъ|-䧅��ľ��DG1�	���w�/���qΓ��%�� �A/��?����I��7��̗³�=���y9FNj�՗@�<Ө�� =�bgђ)	a�(©���
|� ���0�w�L%can�H�Գ��^9�~�
�ƞ�!�'������',����oɽ;���sĞ�b$��d��0�����p溨��.�RϾ,�l���.]:R�?0~���e2��H0@cD�z>�"т�	�t)Be	��É�'iZz� ��YD�6;�rl����K��͎Ӓpyohi97з�f���߷7l}�����x����:(i��)��f�U͙�j���n0�%��pm��J��m2��XOW#�$��_�ʫ��
��ۛh(u����&BI��Pa�İ�TU�?�p�vL�X�x������"&7h����N��x`(-֙�j/OH�/�����v8�,��[��|�o���K�fѠ�w��V\���>�UMA�B���o���M�a~WA�3��ń����g�{�͓l��$S���*�S�*��F�
K�Yl�~G$�t���[n��غ�R� 톽���)��-0e����)v�^��0�2�Ra(��G���P�l�P�q�i;���;=����`��<�m���K�L>����7n���C��R��� 4�A��G�n��g�j�)u4F������&��^t���g���(�y����p<2b;��u�@Q�7o<�"h8ȏ� ����F�p+6�omO:N4�9}�[T���̐([��S"9D"=��Z�>��k��5�}x!x=8�h��c�_HݢGv��t n|�l9�@,�9�C�,^�C��2ʖ<��������p��������Noa�:s��ed�?�x(9C�)�~$xi9�U��Yt��F�v�c>%+r������?)�J`N��6��U��h��~6%�cj{|
q�h�<C]"�����^7R�nsA�"��b��W�#Iq�WX���0��lI�j��9���g+�����IH���eϢ����l��m�����M��,Ӛ��N�&d�K�M/���L�� L�֨��s�y�]@+]�0B�+\��}ֹ�d�v��,ֵ��6�5'�>�ch՞̜n�>zsP��Է�e�]�<0�ۋ
�P]؃�Z�2T�)A�!�No����h� M�h�*9���B�qZ��n���O�x\�����/h�
�g�Mp�/Y)���Q��V.��pfx�.��Y�h6�]ږ�����f��#��B�����-��0��O�l'÷���WW��*�|�z5��M��r���SǪ��DcIB'NX�.��?ȇ�M_�^>�z"8�ґ?<E����#�u6�k;j�(�ڧ���Z��ɴݼRi��]���(�G��ir0HR4�g�gd#���d���9�T0�;˧�n40���H-�/��=:�44��`���L �����'�iP�?
Cڷ�]|w]I~L����5��Ay��띀,!�	����Wt��Ôi���TH)I�(���2��o�]�{dS�H��:DQ��a�%_�D�9��"0�m"�>Y����)�k��U��ڍolB��y��R ݥ"f���j��_�'�D��7Q=*H��9�gb�%�U0�VJKӿ@1�r+i�u��AlJ�9�+-#❖r$�r�@�U�(S$P�r�;�E�D(8��X��nD��A7�����j9x����Q��*EĚX�eч�H�Iu���U��7���j�&O8Q���Ce8��މp��*��٩6=���N��ϲ�n��g�f����,U�e$�[�m	'�� �65�ߜI\��/@d3���ɭ<���/i$%`u&�E���i9��@R�\�~�F�٠l�3���Y_�2���`�)�-T����ǎ!�Z�!˷�����a�����k�����M���-~�����2eGD��9��#ڕ'�&��d�Oi&qF_d�Κ�uF�\�g�'k,����x2��@�x%���B��Ѣ����#83f`"wR�s�DJ�wF>]�#VMdDK��|��oI�#�Z�9�e0�^<N�ݬ�jsz��[e��{ ����!
�:�Q�V��;�CR�rѸ�K��q������e y�^��|e8/�)|XHu�H'�[����;o�`�� ����KB��@P����aNv.����	��h�9�*uQ���B�P#��(�FUΆk�Y�z��'��h��qOYA��;VI��D��7��<
N����S��?��\3��wCfͭ�0�)K{��Fr<�=����*�>�?���R+���'��4Վ�<��k���'(��Q��[��o;�N��E��{�4���=���S��}A�v�a�y����!ރ5�d�:h�5y�'�P?��j���j̝ʔ|>,���M��P�<��sQ�`/�7[��R��]!H�:���` %�ټ��Q"��_:`�~S_R��.��c�H
��}���R�btQb���Sv ����)Q�#^��{oj$ϯ�7�,b�fd��W�
��C���'u�ݐs��0���UE��"Ҍ�h��������3u��^,���E�����W�Ca߶��
v=��'E�v<�b�fu�4̰�c��ơ�Q��`= �����xS�W#�I�oZd�B��7�O˷7iK ���F���a��w���!��rH�g�i�a�	{��������V[���{�ַ)�����
�����U����k+�m���X�
��W�W�H Y�ҋ}��Ou��n��?i�fّ� ��x�TqM�F�V�����Ky�؈g�Y�$�Q^���s�[�c�(��ET=��Q�.�2�n��&�O�1�;r��_�<����������	A�_�L��v.46�^�{�?p��g�2�L���)Oz��ݗ�B�9� +�h�s�K��7���Od�T�عu�fW�9T��@vV�w��7�����t0�뢡b+_v�=�J�%vFy�B5����Եf��ľUA���k��o�Z9���274K��і'�[�'�]4yg�8����z,]ߋ������#���MZ��)���k�e���P�)DǍ��ޖY8���yQ"@��!O���F�
�KQNP��u�gWo3V��t���N`�"/�J�Qz�ό�&E�5�؂�5r��<��C�?�Hx!��Q~2�l�mQ�C�-�K1�d5g���{yP�����X`5�O������h�=����#�f|���4t�ӧM�ε-��.Ō�J]¿��MDGa�Q`���k�����q_/���KKx�������/ �"��,�ʻ��'d"�w�����M������/Jߖ��0���(���K�_�2���
5&2��,u��\# �ع�+Wm쬵|��A�yW1cDG�#�/[K�
i6��q���v����j}���=��6 "����rԿ����9'Y�-D9���g3��QLd��D��?���X]1F���ʾ�Qu�@��_�1��ֽ���UF��D��/^�U����W�M)�G��=���"=�+Ȕ��FG�%"\�*P6J��������쨊�[}5�K}$�Hi�H6F�*�I����/�R_�!�����G��3p�Ҩ�QU/�R����
i`㓞�o�A͋��G��Q?,y�F��<+5ɤ0-�)���bv�ؖH���(�$d��o�G���0�q�Ib�t
��S3�|c���9>,��q��)�C���^��a̻ܗ�R�g$��ϻ��)1]�5 �ɧ�N���ec__O��iv�oe���T�<\��Oh=�X �� ?�M�w4���c��yA�����r ib&�=�%�Qc0D��X 0I{�zf&IX���`�����_*m�w�<W�x>��Ŵ<LW5τlo���TCe9�dyF����~�a�z��꽃:���@H �F�*4�>?բy�:��&�d��3��y+��C�=��������nMs}V+g;E�Ζ���d�6����`D��a��>��
F��L����	b�/挙�Ap�=�(�(�?Cv6R,p�aw|]BZ.�_��pn k>�`�E��Pkg?1���JN��s[?"hD� M�_|'�""sSM�4����)d��Y�t�1�{�C���?5CdY�虣�ȑ9�	Lney�X"W����9)��b��Z(�6��SH{Yb���"
��7�>��ɀ7���պ1�7�ۧP6��(�;�V�U�y��a$���і;'�%�V�{~���٪w���r)aT���d��\)+R]��0��ܽ�DP�;����0�VF��47ܣv��u�.���d��V��@�i)v^Է��GG_��qVxFw#M��ʎ�<]��!��0�bCB�x��0��̱����r�ۑ�TWp�}�N:���a�Y�e�ˀM����pmf�=�R���Z�J���:q�s2�w�~L�x�d[�h�H�!�_AM�,n��A��ޡ1�/�[�)4������o�ZZ��Z�K65s���I�������$B��/�p�T���|���Ď!
]���O�#�b�aʇ�$׽T��+m_���Swg��v^T�Ǉ{a �����d�c�v���L�I��J���BA����w�6�u���*q����i��sH|���͢r(���8��>?��*�k�B�B��Fg�F����Fl�7[y��P7fO��,��Ϳ�hԊ�m@�D��VD+����7��e,7N��+X��T�W�7:��H�A=��kV��)xz|ϸc�z\��d�}{A:�h�ɽ9�2��=
v0/�¢�(�H���q^
�ެ޹R�l�|�jd�4K+��{�8��ڐ�ęT��>�V��}�@C��bwc#tׂ��Kw؆�d�(5[�#���eM������nM��|�OS&�؄7�%����g�4$C(��Y�`6|�CS���䶵�a91�d�{��%�?sb�N�N:��y)���Pc��6���M�O9�\�J���c��Ot�~�Bsi'di�7�6�����S���ԍ:Z��n�D�D�Y�����sT=f_�t�1A������g��<��
�;�� �{U5l���rvvyњ|Q���!���Þ��V��cԉ�݄��X�I$���ݸ��x��7;;�{<�6�Y:e�p裂"���c�F�]�L#_5��4�  <D��L�׃9�&,�f.쇱��f�
���.%��ۘ�N%�HZ�9ȥ�����\q���h%��^@�N��$,-�����" [�6fG��1�"�8�V͵�L�ɀ��EpU�stʛ=I���.f��Ag��:�	~Nm��ʐ
2� �pƏ�Y#�,��  A"��#K�8�}Q�[����<�ѿuwg@�4�H��u�pru=Y�v���P#T��,��f@��˫��Ok�C�M��� �Lll����C)!�u6�=�:�Ny�c{�`S'y���	֥"~�H甒Q� ���2 ��|���r��R=�� ^V���X<���UX���L�
hg�X�M���ha*i1n��J�YO�$+�6NN�a�Wre�����z�}�#�q ���N��esq1X��״�=贆ԋ�h!�7i�"Q�dP�WX�̄a hn�dT�j�P�����I��"��y�փx4���MO�x��6ɿ�_�i�����X��m�\�W6���מ��~KV����r,M��J�tq7G<�b�7v�
���e���Kڟp��P�XP��Õ��ϭ��G^ߡ����<e�2c�a��=�@�-����|O��ָ(d�%qZC�&*�u�^]�o����X�H���v��_�[_vW���� uy]_�����e�Dm<"�2W��]�C�	&�_0�[Lno�Yԭ	��ъ�����/�}�S�G�����@PP��;�ɓ1�γ0@���`RxQ�doy@���`�=t�0�q�1O��jiV�7u��Y���/JP�$�7aSic���S�s1$79�����wK-�.U	����<�����
ٚ�p���r|�`N0��W��s&���G��D�����D�X+�~Ŕȟ,qi�L̀�޲]�j:�ui�WE3���[�!x�g��������	x'�]@ᆞ�'T�1v�?�)����EdJc.���V����vʽ6}�e7�p�tk�d�����>/bݳ^uWR�.� F�y���ܣER�	D��{��~[�p9�ջC1�'�'�Q9�ꔝ��U-��/��*�AJ���≻��K���4��?�,�`Si����v�"XD+))0������U���׎b9?Kކ�9����"��*�¨�9q����v����8�#f��*�:���ɝ�0��JڢcM@��'����@
�+ܻ٘�ɕߖwr3���.)z��S�����y2O��F2R#`������Y��Ó�a��HP�7J�Y��B��;g��>��Oh��dJp f��q/(L��ߛ �-�:�Z��0xq��s�=�귺��;�b�r��Ԙ*��K��)����i;k�?!b��.��֒T^���z�ieϴ����=DS{��i����f��5T�(7����'���&�.�!��Of����%:]��v��K���D�j�ɜ�<��H�5P�ڽ3�U���͈ ��>�W���uk�GsfߖH��A�|6ʿS"��'����Zy/��)��~��96^b��g'f�ddBpo�nٷ�B��} `�K����H��R4�cU>on���7��GB�ؼ$�H8��1�C�;0Tq�~{OJR̼�������x��4���j264����,����t��n:j�.�qnt(
m���1�������du��pu��'ta[r�� ���6O4ke�	�:�t�L��	�=�����nw�P��Us^������3B4�#[^{�t.���9p@�AGp�ُI,�U�Y8��r�n*���4���6Ќ=�4�+���\>�̢�r�|
�{�8��enx#�D&�x���Ss�
����;quW�'s� n��6I�K�#/�!�S6�Ep� �Y�12�7o�R�Jt�{,��ړ
����f�>'K(X���S����ɨI8���|Ǌ�C��K ���Q#��f�GM��Kx�EB��{R��|&��KA<�����z�l��5*)y|.�n���F
��w��m�l�C�����k�l�L�}gi�ɎO� 1 F��wD=��5;���`B_���g/ȀwH
��Y������FJ��0�s ���ȭ�i��vƿ
��G��	�쁅ZA�<&�:��b_N٥�����:_+y��$�\_5ug��V���0̋�W7t�]Xq[�_)��RzF������ƴ2 ��X)��y�l3��Z���UC�:0��K�<9D=��_4��p.k����G�|R4;՜��Mq��i�TN����"NRD��}A�x�,2��������u�ig�H~P���ßf�0�i��
��x�ď����2<h�.!�����	�*
�RFE"(lZ�X�t����B�z��}�������<����K�ލ����f �"�,�a[)��<�h�!@tk�ѓ�Z^k1(J,g�B�V%����E��鐃y���P�W���ڷgZ�!S�#�ۭ�����*F#����,W	�L,��m�D��w���z�/����v��<p!p���,����k��n���A-�|uP�ri�|�A)n�=3ۈ!�g:����M-8
��aC��5Lg�[�I���{�����1xzӷ��4�E�����g�d8z]C��!5�Tl���=;C����w��4�b=|�IؘP���bR���͉fO;����5{g����W��=�������`P�`nNe����)NkJ�5v�$��p���-�Z��	\���	*.�PxC��&z�q�攘k_���n~K,|��_��v�Qiê{`��T��!a�x+��.��!7��5��T����)p��������yXYϥO�GTͨ��f���s��$�W����� F/��?l�*J�?7G�d�mT�G��(���n��?NO�W�-���$�p�m��j͜c����\@�k�S��_ڵX��+V�����n$���W<�˱��Zs�OP��S_� ���k0n�Ľ�3���dʏPJwNQ>�3�u@H�ac�YZ�Eֹ���/&�y ��s��R��4��>)]�Pyj�����B��".E�թ`-�jZZ�p����s����`	�}�:W�f�g�E�H�u�/=����f[I:��׏�3 SCa=��16�\yx���zƾNa�L���p\
M!1B��B����z=���pU��?���G J�7J;h��C ��}��z	��<q�����
�"�	�FK��8�P�۽}Ӕ�����	�D_!0�����
}W�,3-���҆R�g�Jʐ���ٽl++@N�|�BD�j�5lScX��͸�+��kg-j������BHTnH�;�tf��C*���e�Y����?\�WwS��u�fK�cM_ ��S��.�"9Y��a�� $⟢0���"�6;�����R�C�Nн"KE4��$/%~��w��ě,����n�V#����a�
��4>�N�;|���_���gV!�A,��[���jFŰ.[dq �tD�F����+<0ia�SNW�q�a�1%��[��%�;�[L�Z�����Wu�p1��Q:zX�#�'�������V4�x�B!��)ų՚���e�17�Bл�2j˹�V�|�Bvu�֎���f�'B]nt������#�2}�7�R�b�J{��%�c�R>��mu��y��L����P�d�l,��)��� M����R`�ٌ6��;~�)o���چ��~	l!�|��S�-�~���N v��	]#�5ߙ�AM �5�$�`�Q�cncJ Z��-��$8 ��_��O�\�0-�E�b�#K��R�@~�>�e��SY���i��C�ޤ|�o��$�Ȟ��ˎv�@ǋ��<F��۰��WS���}�E`D�<�� �o9C�i�#7�|kCvǖ(����H��i`�w�yj�'��r@�6�Ǖ7(�����L!dV0*;�A;�&`P}�߃R Y���}�n�[���.���� ��(�h40��'���}*�y'F��|O�%TG��P\��9h~�or{4c�ǰpd-��W
�Ң��'?(��u�p��b�w�=�4�Ȁ��1�L���J� �`�m9��:1xm�܀��T��-��f����?h��.D���8�x��Sq��Q��@��V8#�Q��F��0W�y�+��7��$�=��K#�h�i��s5�U{n�H��&��C;�L���#�X�Y���R�#�\t��@��f�j��0�x0
nw�4�}U�8�����(%*w������R������`��(؉З«	�	qwRA��g�~qJ����VQ��Բ|���z0I}�������_��,m���C��z��.�4��tv�"GWr�#����b��Td9�D�^�M�`�B� �jW%I�(�ʲX���θ(��)�k��W�����3�쵠٦^� �C0��?�B�8@_Z$��s.=I�a+�TrA'�䎝��"��g^��NLS��3/��85�[ٟ��}��ϩ���~�hfL��A",Sw��Tn�@��8������Z�h�R?���Sk؊�d0>��y�5�X��8���k�����P^+�ۋȌDH�Ϟh1~i�Vw���$�������'���/)*��M`�Mc h2κ����B��[�75�m�zp	�n�f\����[��W�q��F	��ߓ�(�eCR���8P��0���T��&��I'��:	\��,���	�*_0��R�	)�Nyi}��=�-?�_sg�k�H"����~&t��g�Z�*��ԫ^,Le�ҿf5���$$��c��ب�@׭n�YGq  %䨙���e3�/}��(ńY����+�Z�F�I��L祇򥄡��hWi�����?aWD䱴������{e�C
z�[�zj�Oq��¢A�����uګi�{�@��j3 .��y�����jTf��C����N�ʠd�v�G��x[O�C�$(G�g�aul9+�������^ �`�F�g�K7Gn�UyD\�ܨ�h����$��� ����~�ޞ�j���"v�U��L�QLݣk(�n0�D�)-��ϵ],��R�U
��ͺ�;�t���������X13x0p�u�q�䴈�)�������
����$J��N��rL�@"�n�%��g~�L�sh��&/��Вi��Q��d���8!.C���ږT��D@I�h�89��9Ҽ[{�+4dF�|�d5� �����C}����øuYP�h��!�8,����L��wJ��`+�^y3'Fn\�w�xU���P}�p��
��0��bv��\<�?���~���h��-��Ԋr�$>M�A�����}N�����]��wܤ֙zi�O*�l�Lp�:��&�'��,���q�T��<�������Si��Β��nf��-7MŅ&�t�+�����/;#:a	th����]�3�c�ց��N��,^���U�Ţ#7�T#�/�N���WBe����3�*-s K��4^�޼!ꕱ�u�Ե9A���GP��9�w2��� 'KW�+����8�?53̉�����������8rCB�h;]/�h8�:I�8��1�=lr��� �QI_KWq�B[e���M�$��0�r�{��侧U��)���З��g_T[�r#�c�2��Ĉ�.HL^2n;�].ڥ�"��+0�5hw���0e���C1�� �!�3ВC(v� Z��l�X1?W�	�r4eu�Պ4��1P �����a���S��ef=L��?�(��[�P9�����'�a
�ؒ���EW�>n|m
E�c��+|ȍ �������d��R*S��b-�o�B$��Lt����A����U����fZ#�Ė��t;�I�
�?H�i�b��z�p<����$�w�!$	�e4j�.��џI��u4��iI)ղ9d���G��dJ�@'��ƶ^��k�[��C?TO�S��OT���T�^�X��rxR�����T�[zB��Ŧ�:��+D�4��u�	���琂>	��D���u%�JYva�r;��D���l`HeŲ�H����*�q��[�X�?0��-����A��&�]�Ǯv�\�'�~�u:��3��(�.������f�`�d�Ǿ�E�m�վ
܀_;�)�c�nZ���-�ى��8��0�]�<��mw/���mi\Rqƭ<�{�&�8v�5i�l3�TşS�>7�.W�3闞��>���p�5.ř[ht�u�J3C%��`����9��'m�S����:� ĩ����<l�L��l���k~4@�]�p~�	��eI0�	��<u�M9����7��q(�`�ڦd4��~J�����2�g���F��/y�D�=�P�z���(n)m8���&*�8��5��~��շh��k������P`���[w�5b����)G�͙��8�Z(Ho�5 
� ��i��*�̡T�.3SJ�eIi8lwt�lpPn�Ƙ�%򷼑�����^�+:/"/���t<
��:5��t��x�<$�p��U���H=D~�ɽ���-���+�'-(�q�w��L���ȉ�t	%���z�E�M�N�3�>��`w�����$���4���l� ^�mNv���3T�m���*(�`��Oо�#�'Ƿ��wM��v��K�0�)Hr/b�S3��B���G7XPFx�k{,��eզ����C.��0���p���=�4�D��N�͘�=�י�H�`���V6�8��SZ�3��9��ϑ��!���D�2�.�k�G�0�������2D���%]�J��[xR���N��٪��+0��'�=W�ٵ!!kP߀2Q~�b`b��	Kc�����Y=�Xk��<�t���ؓ�ۉB�%�w��hᅽw-jˬ�F��5=p1;j�h�\�e���I��Yka�/��{`��(�[2b֚���cvYs7��ԟ�	DXO�zLw���p�v���b���>�2=��a�5�
�bQ��Oym�GA2�y��pk��.�f���\�ɓxi�b����(��S�+> 	c�X�8(�c~@��
�?ݠ�d��D>�`��4���!��V�����2UD6�Ė"�
q�b �*ϳM�?h��������q������AG�W�/�t�/j=���h�y3�@��D�y�S��]S$��	�x�@"��� �9�)D�:m��1�T�����@*��R�
��ud������B��̂�y.̝S�Q����A���b3��A�yNAťEhx6���-z_�
��GB�cy-�D�r'��y�ţ$h{�G��c�6o�YԈ��`~��h��4hv��*yO9�2� ��ϙWqW~gn� W8���ki,
��EK�Ll�}��`��^|&>�a!a���Y�|�)%)6��F��U��J�Q�5�:u�oI#���؄�7梭<Z�VF�њr��b��$��bze�Q�[���P R ֋��!�jj4���Yx�s?>�ҊZ��0`wF��c�A��%���i�.��z�ļÎ��U�6���7�G����3>C� ������Pԝ�c���.#)��~�����V�:vi�������^��h7�n�G��1fC�ɐ����h �դ.�]��������
	���q�!����(<�J���[J2�o��vnc��[
��v��E���6������{S1EQ��o~\#
�<YJ0��H��Nt�S������ݦ�`�5M��+�x;�8ah�͠�p�MK..���ٿ7�\H�wZ���9��w7�U˹+��{�^U�d�b��s2���엨�y1�����?�.�e{�:��PT�H��(�l�r�_�[��ik���Fd��%c���ͨvp@���â��$��uR48�'2ZRA��l^B��<�ƞ��Z��׾�Q�c���sT�W�'G=]���>���ɨ��Ł��g�l5����*T�S�150;�]��'+a�lh6:����L�*_����dTp1�XB�F��v?�6~�"NB�6�q��z��	���-/��2奼Q�X��$�%���Ę(?��Tς\ŬW ���,i�yOҞ�C��[��ji�[t�������f��ND׀HG���1�,^ �M�y�$�w���x�^-O��.�m:�]|�ܓE���jh�~>��H��0��l��U+'^�SԴ���}]�8x��4sMLf��C���5v�e�D~���������>Q6��������\�Y>x�Ϳ�����Gh�@�8��B`�m���&�L�^�G�R��	0(FR��k���|!��L��H�_6�b���Lh�����nd{�����sԼ�z_�,PL
bzS������(���,�w�M5�|>�٢Ն�J����#Kp�#Bxh⌿���ځ�6��.���%P��<qtec�u�e-��'�'��I��*mO�j޲s�XhY�������z��ײ�9�,�%�L���t�f��>��Ǖ
�8��	an�]�=�g�lU��`��y��.�w���<��w(�![�v�D�_�YJ& 
V�ò`����{9�p���)�rT�v�Lr;��`���*�+:��H�)�#����E ��)�Yn��1���m�j�C��1��N��5��B����l����P����������U������]`�O�� ��{]�Ƥd�\���:qnPeS�T��Cqk�����=��l�����G��Y����\O�ۆ �r�'aȷ4�҃������k��آ	9�>��u�Jx�e䢰����$�2}ߨ�n�p����?���ٳ5NKɃj����]S�&Y(X:�i�oٿF�jK�Z�3�Wze$d����G�Y$��1Mxl������5��<�a�����n���<���r/MqHxr֌����a=�����[���_:}��N	:\��ʱn�r%L�`������]G�3������G��̔Pcs����5�K�7yK&V��_�g�:k<S���C �
7��A�����d����c4���"1�11Ԙ4��0�b����8�dE��#��|�t
-�L�}����Ƥ�a�U��D0���;�ͻ>g6��8���s��E�WE��*7#�@�����p5-7��ҭɔ��!�,��x�/����k�:�jRi}$$'V~\�s�q�a�)�L��k��'��mo-l�G�u�m�5��nM ���";�{�#OZ��mWT������҅iS�3B�-[`8M�-mt���	�>�,��R��pj缰ݼ'?�w��7�î]�xz.pd{OR �]Bd���ٵ�k��%�{����J
�ɚ�TP�r�)I�#&�":$R4����E ɡ Ӳ��]��KR�}3�'0l��Xc��:E�^e)���M p��RM`_F�=
�	�(�}��*�T>Ǩn��)w~L��A��qb�.d~�ײn$���A1z���YEc�����ǧ/��'4��Ufpg���A-\�DŶ]��LM7�̺�C W�'��j��J���]l������9�6j����6�]�6��b��$��+Bí�d��Զ�Ԇ*�
5~�>�JBi�$�<�iho{7�]����Guv暥�8f]%��u	�1�m�͆����4>�l1n%\y���
E�G�\���si��p1.�c��\�@�r�Z�B򘮹��NK�B��Ƌ\O�a���� �?�o�	V��ߣ��ڬxH���@�����5�n�3�
nW��ڧ^�ߖrǎy����K�fo~]6r��Ҹ��l��N� �-���[ �8AŐd^=c ���i�D�~ %�FP����CA�7J3�m$�9Ȁ>\�dE�d��Sv �L��Wf�R��2;5q��X`v��%BW��1G�ezl����67��x*�,wYk�3:��ֈO0C��(y.����Ũ���t�3Xi���|Z�V�Qh"
8�#'�E���b*�lh3����Vg^�0&#�0�Dm�L�R�+R��u��W)��X�n2�g��i���AY�!���E:t��52�/]_�����Q	\�[�hn"Z/M�8��DY`g�|������s�Q4pH
�|�
!�9�?m��iM�Bw��9N+TM��֔⏕�á��kd^�K�c+�)�m!Af�T>S�[R��8Bd������gA>���.2T� ��6n�+��j㳺��fʪ�¨��z�f"q���A��B,l����s�'�$�cZ�L������[1:}�l���^:���
98���k~)�ڝ�;����R�8�:�3�� hp$��(���W�WVT
����əl�֙t�!��Fߞ���$8��w�ׁ+¾7�HB���"� {�9G\.��D"K�ڮ,�O"��EY��|q��3i��\��*oz�ŷ��,_Pk-9<���/�qf�Wb�9O�L�)�U�!�M�z$�&"�}`Y�?S��P褭=s}�O�C�QQ��le"[^�)L4����cx��~� L��), �u 
Xҷ�1��_u���J�>�;�5���Py����!���AQ����o(�g�ݰ��'�˄?j̥�NN��A=�j����-��g����HO>P����j�ץ?��` ��(�g�! -���4�5	3.㨎�5G�l�+��E"�7�j�StlOfr��i�=��rUm������e�x6���Uߍ�'�u�Ծ�v�*A���MU��Y��/��.�N�*�O��q�>Ek��������Pȗ��j!B��O�E���}��͛7�h���V�]a�:M8�M�$2��u���l��b�3�}w��of���6�r���)[JjpΏ�6���� O��Z�'��'��]�������A�Ϲ���.J�E!�����iv��T& ޽��X���i̗c��u��S(���>���Y�~vOa�Ԟ|��K�ꓣ����$� �np��rU�B>��"���9���҉a�e&hO%�M�U���Q��f�I��3Y�ܧ��5huc^�?mv3��L���"��[�+.Qc2�� ��Ϸ��J���C�J�՝%���֙�E�]�湷~����Z֪[O̔�o4��.��=)����}M);_�p�v-9�z��1�2�x�d�7)_�Y	�iٚ}�Guͧ�a��jKA!�ΰ4��G�Fi���nd��Ȱ�}�O%�6p֖��!��o��2�����`x�Dײ�&)��s���GU�����D괾�4�D29��j�|��	�;��;O�
�3����~����[�͖L�� ߠ� O���1rcH�����w=M��~�D[g´���4Ś4���1�	�-CHW��A�Sׄ���V@oK[�i�[���]c���sĈ�J��ď~�Q?Y�3	0LU�GC?�/V�4ª�!�B�����_C���H@���7UQN�ʭ��i�A�~$�%:��J�������t�?�� ���L���8�^ӼGin���@~�@\#�/��r������;Q���xEK[T;:/�	!AK��L�c7���)���'u�[�zT��"N�{x��8o����t����Z�OԽ��cs�5f�W���9ڕ6�1�O���.��\a���E.�h�:Ӏ��(9�pHFxH�n<S��v;��B(*먡��cUj!pb�z"t(��}�^��3�vzG�Nrs�J(�������[�n6���=�@(;�P��fS�1��i�{�L%v�>ohى�1�_������Τ+�����q@�Т��5]�R����"��}�^��U0�\�'2~�ӳ��=[�ery�������,ϣ5���wO6.�8Y�,(av���{�I�wpu�'epo�o#l?�7�``fk�������0A��tB��e��P���ǳ��T��jP	��Z���~U@��^n:R�{V$b֖���W
 0�t��O0D��ɸ !ڢL�9�x��ϱJ�5���w<4w���!��AHK��8��V�p��H��kF���v�-��?��ձ�P,K^d�V��N����̪�+3,���/�C�z� �����.J�$����x��R��I��+�-���Ѧ����w�{}��-�.k�hX};�Ͼi��b"m����s\����b�d�BS|����a�Q&��f��I��uy�%!5ɮm�I��u
j�����3_;�+��z� b���[|]קX@�d|�^���\�^W��>�Rڊ�����l��ο�
"��d�IW@�T*g"с�����F<��\�7�G4&.��>���L��\��\\]��/m3��T;���g�A�Y���۝���/�u�݂H�_��l�N}�U�6D$�By��s��t�����9)ЊU�����p�[��q���?�L�\R��bݓ&<g6�3=�Β�B�X�Mm�)�sC�^�w��D�x�Ĵ7�ݚ�0���*��р@4LNGlw����_������R��;��6n��W�t������q����LF�)��7z����bp/|�j��|����R����X���k����O�ꃫ���|�yC�P\�	0�k�zʪ���b-i�rƾEܵq�"�hC�^�yk1���~]aΦ��BH��5v>F���T���M��?ey����P���［'�r��6��*�Jٽ=��}( �(�T��91G�WyI���Ղ%����ئ)!`	2�t� ����U& 7�=O�îE����2�1�Lb�q���C��D��n�F(i�JJ)PtJj�ɐSZ/x.��JݓXj\ĺ�|Y}���W�0���i�p��\d6>ӎ#��6��%ˡrY[*��X$���@3�òO���A�
$����An�����N��G���;�����)�l�@&��I�THzP_UJ��r$*����[c�k��?$�yJE��B��Un}�]~�B ��w��,��]o�_>pX��!�w�A\��=��d�aZ`���T�F�`�p����f�]�|����V����u���윅DEd��Ҥ�:����J�U����c<ůq�<�����9Jt�7��dSG�(ʪf�"���7�/��QFf Ň���"ʡAwcgY��?�M�>,v��#k$A9Qfm�1�L �)y4 �M4&���;��Y��S��-�E�I�R
�a��%�o�@PsE,��3�I��X��G<�m�K6�s��kX.��l�f��<xv9\��_��ӧ�:l���-?�O�3=�P^�}�]���?�щ����P�u�/��+x0O
���ח�����/�)�yBl[���7���ß	�E9���LJ�{�&������7�\}��r�&u���(��Sp�� Y��}f���"��z8��� �g�75w��W��Z:�wN�س�񸐵<Cܛ���c�L�k@*C��6JĦ]��+N�0!T&f�GC���ho��y
�*X��;������&�/ޤv�C#�����[2�gH�Pl>��\Kl��R��WP�(6��>X;�}~������N�y��"*�/�2�� E��b�,\�?L�����rs���̈/��^��a�)	�5�6�Ŋ�һ�K��l��l���u�q��2����c$%��zs���X'P�|�ugv�x���:Dw)����I ��c� w��h���ↂu��uߵ�\�������I^Ws��E�Rژ��xA2��稳�&x�k����D3��>���n��u�3}�n�������yy���1^5Y~m7|���Z(��� ����5�L	�[-WE���ͫg-�˘�ph���(q��Ѻ*ζ�\�<���JH��˕ڭ�wK_�|SJ[ )�1��{������SJ�����$c���/٨�GG�b���\c�k�q�Ňֶ,���|�ym[��5�YiG-�aZ�qF������q��d�цg�ܕ(�{��c�/�9k,ªT�=�M�Hl���q�ZRǕ#����� a����f��iv�B�6�/�����Y�6��[��a��Hm?\���nL����n�Xw�bX��1����1�`��N��W�WBO��O=��2��>tˈ/��"�@Վn��>�v�%���u[%�6��w���?cY�U/�
)qM����K\G9U����W3����J�8��8�`�!@����yotd�p�ǒd4��'��c�'���u����B��.Nv��ͧ�+��D�ڐ @)��i(1��"�r�_��?7�j�z-����?1�%K*�e<����.ќ�98d@Xȃ��]=�8���U��35q��}K�:�H�~�ag7��A ��*|U�M����LW�c���y8M����L0�ݟ5�U��+U57ؼ���@��)��y{��P�R�)l��X�������>fP	��yg����/��$D-�#y��im���C�f��y�;���R�l]�?�AG�d���\��������FV�g���W������I���>U}��w�b��I��
mW��S6�c_�һQPq��p%zV����Il��cddM\�JCR�v+��e��	�z�A�+#��+V���]@�������j�1/p��'��r�g�{�=]�q�����#�L��^�=� O8��)�7���(p�s����_e��ț�x�a'i��'j���y4#�i��I��[6I�:*o�ޣ�~^����,���.�u���_M#|s1'�7�!w��b�nK	���D��\`eN!�B0�ߑ�N]���6i�x �b��� |�c-7t�U*�M@/b�}{K�N�Md�,V���&��_�9���;?r�G a��Y����IN*�]�7��� �s%n�h_$��}�pdGE�1�A}&&,�B�.��?�c���S2�E�R���4�*��Zѭc)u�6�vW�ڼ�bR]%jg{K��V�,��`�&�*�u��Ɏ_�6}�NEϧy�4���t�t�C~�:8�ᄸ���à=˚vn��`i4?)\��̴��҂��R��Д�/a{�n��8���5(ŭl�~�祿��|�w*c��7�k�cU���ܘ�\TĆ���Z�d�a����\6�m��r:�[���4���@���]>��jݸ�J0��edH[k}Z������z��>y嵤����l@����a*J�)�k��8����Ӵ�zt�P*P��w�B�����E��g��U����\(Z(���j��K.&��Q�����+�:})�Rm����|D�̷�i���gH�*�O�+���|�YT�!��. �:W�!pѨL��7�7��֢�x�B�ݹB   ��e�I	]��}�B�bv�h_i�c�'�4��IK�cOk%�/v鉵Lc|U�N����������Z��s�&(�zN`{_��f�~d���8C;I5;�<ɂXe��{~#�1� f�d�"{�U#��=�k�E`�~dɴ��	�h�m��
�6D>�W$�cGz���:��iT�@x� �Ø����	6s���V�5���i�H*�yY�]�����E3��O�>k ��HdCEN��d8Ʒ���~+;�c�w����%�
/0�©����9�@q Z);0m3e,N��@���'H����^�
+�8ت>�����`�����X����76\f�q�b���n�����m����ڞ@��@�V�6V��z����,��0�����e�ᴼ<7��x�tC��W�;u������`4�z~vX_���gx�٧D١s  iؚ��89�>mJ�f���M�Yi���b��Ef�\JL��؏R����xs����u~�`umh�ϑ"���Z�nL0�� �Dn.=+F;�j8�wC7i�}�V!u>��I:9����p��v����E�zL��ݟ}!M�:<\��;qP�J�d�R���W��
S��K[��]NP����lOm
�6��W#�O�{�$.>2lm�շsY�½fQ�Dt�v�Lo�F�<���{��1+����	1�V`
�JB[Py1�k��p '�GF�h��ʆ��G]x��-�L�CX�_A���|D}�x�h|��Kz�ؾ���L����&���@%K���K��`�%H�iY��ME��\|VD���c���^wUg��3f��x�c5�*\�ꈄP��q�)��(+���k�G�
p%$W�j+�����O��d_C�P��qp/�"�qd�q\棌,���20�*e�O����P#���٦���}E�Rolr�$��O�}l0K���?�����6:W�ɋ,�&�b&=�%�i&�/P�����ɢ�e��*���y��a���t���#������۾�5OFŇ�Es��}�C��K�ɸ���5���&�+�
Ey��śy܂G��f��cckK<<9$�Q�ű�]���Z\��0U2���y��l�$1�j�đ�R���_�D^������o��H׌��u�H��j�[>buՃC	��(�|�~!s�0���ݧ��M�7@�4X�}�>��������c4NS�����x�B\��/
f��~��*v�Q��ʵ���Ԑp�f����Z
g�3����0#�"&6o��M�]�1�O�U��..� G�c��T�!�ٍ����[��M�a�Aj�ZW�H���s:�5U����ids��6�16�֩��U�-(�3e %)�ۧr�@y�&�y�*c��!�� ��
2s\�M�֏z�$�x5�[�@%F���-�]M���	qͰ��|&�2���3RȦ���5*��b�5������l�>�6e�S�F���o)w-h�]�B��'��D�l��������ވ?�5S<�heezBo��~�͜���ѹ���*�(b��P������IMum:z�����]܁�͚tg��ÀI��Wt�&�����G�N.�q��;�hk��A@��6�\�����ܗ-q��3\5I[C���3�����0A�{3�x~���ϚG�G�t�ۺ:�ORS��H�lSCLl���)��F�|�4c"�GVl�[����/�ށ��� A:�"A�T�c/aZ	��t�i��s�}>�_6ԭ� �6�v}�^5�($s%�p)���GA��cwl�5����Y�{�$� ��Siזx�?~՝7�O*k��z�c��16�1����k��5R.�'�� ��-j�x �yQٕ{�	�٦�A`����w'� Lt]���B��!�N��JSB�X��^�t+Q����H\�G��p�A첪88���^�d�m(��/&�Q�:9���"] ~8����كز֨U�z�����e�h��|i �����c�13.Q3�Q���8��dAC�KG��x@j�2-��o랱�����/K%�@Ҥs{���v�a�0ڎ���L�,����Z{/��0�1�x��<l���]Q��˭��)����a#�.:�j)%���8� �~׵�>��rV	�c7�vRN/:R�}��h|��������P�o5��$^�!y��.큞���w= -�x�,�����;�+^ke������ ٯ�I��xڻ��H���K�9MXæx��19iY��?z��W�|tv�k�`�I3/J�L�����6��7��1�A�reR��'�}c�����X�n9&��dj߆�+�J�r�=n�� X� ps4�qף�����y�h���x��e��#D�L�4*L���eϻ��-:ꗝ�n{�r���rӈ�X�C}+ <N���=�X�d�"�%d��dΉ��hl����3aW%d�G��݀�E=e(Y�D�Hm*�d���׋+��N
(���oT3��DK���Ԯk6�c�؈�r3�}n�Q=�Ism�1���ҿyMn���X����:�8�2�]���G��5i�����[?�/�$ʏ�t��af*�Ed��+�����f��5�i�2��_ ��4��@D�T{]>>!��<���NQ��Y��Nq�AH�L���2j^��g]<�ꊀ�Ǵ��ra�(�����.E_��0��Ȳ��G(G>���5��$��镏۲C�R$���N���d���eu���9?s��r�_C�^����𺳙{�
}JͶ������vӨ)�ktps�ub��D#dc
0�kC.��E�v��}������Zh����5b�+���D���y u�a��
*$�4/�&G�i�H�Պ�z���̩jB�L�I�Z�PlJ��G��'���g�zc���e%�e|���6ԟuQBd�y�Y$@��	.y0@�8�T�t�s�9�*U���� ft�Ϡ�`L<A.�\��ia͞�3�t8���0��a��K�8�Z8V'F>0�G��V*N[��+�}I {�&���8 �hpY��^%����e�]<R�_	�ر�&|�u�PΒ���{���ޅ�[����}��F�h��a+zp�<��t|%�H�ϵ���p���<��{���e���G�0&�m�X�_w��	Ұ(��k��w�����`�F7�
��/ƹ�鿚n<�wg��lõ�b����:���tF�5���2���$s�p0��J�Z�t��k���Dw����QQ�*�Чq��
� xi��uYX-��!�K3������a�SL�"��@Bn�����z��;Nn�[��֌*ID��d�M�����\�-ή0��I��8:Т�l��'�K���4���ķ�y��ZE�/6��Q�0�Y��¸c*�N�u[z��(�4*0�+��I�%HG������V5��3��0�A���>�
=�'�➆�F �j1�x�ڧ��������Vw�o����Y]���q4|p���W�6��·���(!h�����ʾIF[IQ>
?������������2�7P���c�JUj�Y�V�Q@�AC��A���PX�1��H��o����ۮ<��c[c�7]�l�EԖ���R���B.7m��{�X�礊����Ҽ�(^S�`�O	R�@K3"��d{��?��X���Za�
a?��"����lk��c'�ܼ8������ޤ2#�_�k�g�!pk���a���|��5S��\22���xW�'���#�3�;"�G����������2�T�O��( �\˔��#����%����^�=o�@ʇ��[�Ft��v}7�ǋN߀�\Z�}W�es5v���������\.�n�O�V5�*�y �f�t�|��Q��=ge�Ȭ��׎b��Gz�w%�2�u�`�c�q鯖�m�� n��Fy���*�T�hyV��ű��2����hW���fwJ@;&S�'����*���}we,�RTXp��A��eTB��4���q�(��w3%wޙ�Ɽ�@0��}����|b�G��2��+�`O�C�CM�A���mo��U�
V,�f^e\�uH��$�1�쉗�tݨ5������bN��L�zV�!X�d'},Bc����#GEK���\r�����6��Bv�j)k3*G����<�}_˝��79׬��/�j��,t�h���<N�O��<f�kU��P��9�)���ʐ�Te!h���m�M������Q4��g���_q��U{�r��u�e�l�c��z�ϱ���DI�_m�����{(-��7����"wY�����.hK���kva�`9���椁�����9��k<6�tY㺹裰��`n���ܩ��������H���f;���(��%��QN;7^|��糤͝�k	o�������O
_8�Vژ������^�?<|�/�jim�� J@&o�Ql;��O~���O�&��d|$�O�����ɓ�}8>r��ᚰŉ7�>��N�m��_m�l+K����?���nm���`������\0#$�yu��)b�(�Ƶ��m�s7�;j�>��	�Ȣ�Z�]7$��OT����B[��l���.��-�T��.[[�ao^[A�"(����4�Rԍ�f�4�ƭN����r����:���(��78ܖ�\P��3+k�b�>o�6��f\�y�q�k_�%V�X����r�m�!U�\6F. 81�-8��آ�A���T����p7�{Z���ܠ�!iA:H�����ձ<���E������'��r��fT��o���B)�P���^�f�~M1A���0���ü�;>�C@�.�	��~յ�)��ְ٫�X��T�g������6У�,8xKo$�ɾW԰	�m�|�#>���	j�D���%W���s�;4Q�j�)E��E�6Bs5�n�K�0$�x�������k��]fBbKS����Z�&���ra����l� ���h��L��:4���"����.��Aj<ܦ���笹
�aݬW�����D_:��?*`74�:/r��k�
�(J]Y��To���cc
���AD����"<ًrv��a���A�� QR�B�B�&�$%gn>� 50����da�8�3ڱ�j���%'ɝ��̆�} ��t���C%Y��LE�V_E,
�����If��	�>������v+2�7��� PRdl���>�H�c�hw����G��TH�7Z5�',g�W�%�1�=�w�͇��t
�E��⺥[ހ���t�[9̪%8�=kE�8�)S@;��&8f(_��J���cKur���O,J�UA9�FNO�Q?�w�dbv*�śs��뜐���Ua�~Pi
�L�&�jxZk^���MYU�_�&ӇrUrR?e��s���Tj�DH �@F�F�3�n	�Ճ�'�.�*�2��% C9���<�;��h5$�B1�#ƥ#Y�{��O4�r�qr����]����m�m^%��赟sG_ropD�ϡ(�����[qVQq�U�4%� G .�jz���l~����o��@T�kk�\B@}���1<M�kR�LH��2Ϊ�?�䓆�.=�0SVa�qs��Q"�a6�*����N�T�/^�]��u���A�a��M�åx�
����Lѹ�P0��!��=|���3i���P��f�>�5��|"& ��"�=��;��3	)�,�cA����F�$�+)���������	���Aw��5:ȉ�|c]T�܃~K\cW-�f�/2&��]h��Qg�!DLiɰ;�>��zX���b�7%�ßX�*�}5c��f-0���������̱���lc^9OX�����(2���\xǅ��2�TUQY�_�+b dmF�v��@͝%2P�V�=���~�74��I�r7�	+��+N�<���|�������ؒ7�����*��#Oi����<����U��3O�Y7I�$��(kA���R��K�i�L�����+�@��S�J��/�Ȋ����;l��~��]1_8˨r|D�%��-(�*��O���F�S0�q�	Nu�4|�1��M�4�|<���Aw��>p�)$�e���7�'t]�<(�RH-���/F�̑FL�$+�{M���opNl͔h�*AR�QV�7�
�a�4s�7p	d�PRԅ��WF����r��Y�����	~N�����>�[�2�Jˡ�C���Z^x]�k��\^Y��}+g;L�'Ln&h,��v��V =qoAb�^s܊a��b�<UE�'ex�d�Gc�\�m�t#O}
��e��?�E�FSu�j�NʟY3l�"���4w�'� Z2e��./@5ބ�����;����(�5�q���᝾�Տ��S��۩p�#e1�]�
��d�Xw����-
��c�J���<;y����#H�oN����Yk�/��.	\���#R��<y��7��`v�^�u���<[���#�jQ��Z�1�,���M�ovv��������x�P�V����P��WZ���<��˛Bo�E	��zg�f|G�ֶ�C�|�_�N��H�RS�v�U-�9���0`�����p4��U%�W�sn:Gn���g���-�:"��s�K��nB�ٝ�>3d�lJ�N�;
U���6��.�aMBp�7����R�[l�vG0|��ec��wC�肩�}��ܰf�=�ϓR����.D< �k�	(���/�ƃ����IZ�i3G��ݥ�i�'i��	>y��P'�B�����3|ID)0AH#�-����V8�m!Ļ*�2���z�7��c�:8��g{}L��.�[�V�B�VVUL����f^����x�F5ޞzp�|��F�3Hz���X�k��.�O:N5��%�����K�ݨ=i�L���0m��)y�Jg�F`"��
��)�dhd�'1��T�,bі�pX�����hu��"Fv[����ه��O��.7�p��Ł�0Eҍ��R҃�T{Y��ց;�c�O/�DO��OarK�{5�L(3�����U��:��Ύ��l�����q�=}�6#��ehk�^��(�$=��Z ��+̓�ެ뀉}D>��Y�6�֖�WG��g���ݦ���M�^Þ��[A{�U�k-��g����ڰg�)�K\A���J��>]aWT;-��񖗄�A��^)2$Dt���b��~J�h��!��J��r;�K�n��i�)��b�����A���W��`S7{�/���2��pж�S<"nĹc.1D�N͡�I�1�]	���i�5e��87�W���ڂÑ���]ob�����8���'��2��D�(S��M��ݮ���X��j�<V#�D��1��2ʎ$�b-]����9���/�������G��5��Bb҆�����M"\4X��
阂٠���x�?8��1��>��i�;6��K��MF�M�wW\����_��Km1��>�W�5��!�x� GǇF|��ݏ�[>�-��j{��SM�����ׁDԽ�	O+)H_����-}o�"Ed���%:Y�;�J_�"C�I����^A��a���C�j�O"�qizP�������񿉍�\h&^�� =��ҳlr׼(2���0O�u��?���s�"p����ίFb�,k��~Ti�bۯ2|qE�5:��|;7��)��.i�ю|ݨ�9Jx�Ӊ�/
^ȿ�j�9���:��ĉ�.L��dvZ⦕�F����5��O��RްW��"jUedC��w��{+=7�UmAuy@�$�G�Y�cBo��Mp�@�<�%3�&yjE�QFF�za*F�	�_4otI��['|�6��D�����E�1(,�#���`�S�[�).��%�Q�H1���B���H;<'_��_-��aa��a�@kצܢ��{>Ǆz]�9�� �"��[���������aƸ�����x��՚��{���f�+#!g���n�e��PLo.l!�_�u�`��i�4�(L�Ӏ=�ǈ��$g����[�M��B�\Q��5�Yч#��Bb47_��:�(�ë�;�Lo�[H�4�B�#h%0#5�v[�k,gF�Jh9�V�0�c�E��aP���e�C�'��}�˵��lU�+a��6�v�p�썮W�Q�E<�i����7� ��R�)�m���5W�K���=fh���8�S�<�i�m惨;7�0�ė���@�!�jOX�<�A�ݚg�PLRv�]e\��*����PI�����EطH)͔�MS��ڬQ���k�j���~�[|�_uc=�T�� �r�mh6���LUc*	�r����@�g^�ٜ���[��~��S��&ֻGK��cO�X$���{�{,?�K~�|O3^"���Ƶ<Hj�Co��cV�]�-�|3�ms�'!���e`s�0�`�O9�]���1/*[3��LH�k,��"߸�>}���H��{���L��ӷYӫ�&B(�E�{w������O��D�zHJSR�}�:��g*�C!��Q��/�u��5��X��Q��_�ߍ4�7Ob�7�k?n�na�f�y֚��jnZ����K�Oy�DX%9�6OL�L�|���r��&3p�WʠxH������
`�Q�R%Y8|;��&�ZZ�椷�rޖ��0���TE��0�K�_�.-�0r�P���Ikm�@��+���O�76�h��;qZ�zk!��R�K:66�����#���>��Eu����@M>�db�Oi>�ԛ�`Q��/���{{!�q��dru4BrĒ�x���ۇ��YQZZ��p- �H5rf�E����mp���	��ZL��&:
#'j[��J�y�7['h~�S,��Zlk�n�P
�"��U�&���<��j�� ������/d�m�d�ǡ5���!|Y���҅��%�(�+�A��P}�IVdf��w��.�3Q�%�ڃ8���;?l�?�0�l�/�ʯ�Ʃ�Q]B��!��5�"z=����{�cV�v�^>V�\�æ�2[�
l��,�ń����,;m����LJ�kxx�������7m�Եա���69��/�9�J�X�O�Ĕ<f���f��L��N���}�駪���j���
�E|1
v_,(���$~JvJ� �?�;;�f ��#�~��X�-ξ�6�xMί����n���h[pְ�@"#zEb}�(��
	Ja��ލ���-P�Ԡ���7�|��?�~��L"�)�Z�ך���&�,���j�*8ؗ�Ǚq�Ꝁ1��}�d){��w`3�7�����Hs�9� V���_(����܎��?[(���|�X����:�&��lb�&�X�k/!����%�(y)}�DP#�)�@v�
v9-N�ű!����� r�J�l����ɱ�fVC���ծ`����"ŋ�
���>ZR�Z��~s���C�g���/�����(u1�GQ���}O��â�ɳy���r_S23��4�2f��S�)����,��� �):�s���E�!I�23#f��<�|P����t�{:�Y���9*���%���`�s(ǖ�j
��_Nݤ;�aqR�-0��*���ތ��cy�o�z���Ⱥ�"��&�r��=�K?�/!���>�Eױ;
�G��v����Y�]tt�$��W�4��j7@���;ˏ|�SzƉ���nd&z�lmLS����zuH�lZ_�9n+��֭������^��ġU�K`b��mx�,;�@F�9��}Uw��JrF�h}��W��*�Dx���MԿ,�r'Bm%�o!gы���E2p�"�"���	AR�4�S�!S�������G;=��Bԇ ����g|� ��9B��eD��fW_kBWjgm���9��q���a�=z��n�xD���!b��������_[��휳�~>��'��nʌi� �̻��Ґ �ڛ�dA?#��T�Bm<O��(��ϘBu>+����-Q˙@��FQӃ�u+�b���th�+F4\YUrz7q��hx�u�/f�h"�b-S.ʟ�t�<����=���7<F���XJ�C�ϒ%�f�y��K����N���>R�޿Prbl��aK��Kho�.��}ಘ���Iʢ< �XkX��x8�/��2��aiFl���GY�y�<'��u��oj��M�T�A��}Ad�L���,;�q׶� �Zb�l�HSj��*q\��MUJ�FMY�|Q^1*[��T[~��:ή��>��>�D�Bu�$Mb�7�g�ͤ�'T5���&UiC����nZ�_����W!���%��q]��� �p_W]�^Sҏ{���[�c?-sK�h{�Y{H��~�����`+o���x�"��I�e��`���n�X�-��]�P���9���ڷ����0�`�~�W!�PL.D��&�r�G���[Ʊ��`F@����&y�P�ѐ�UP�s�P��;.L�W�&����إS�-9Y�<�κF�~T85��&0�3G-��>�� V C��f �*T�8��[��&Ng���=H���Is9h���f�D��1��-�R�'�������WW�Q�Z�zy�Ԫ_}���l#]�%rԛL� ՞Tx��Y����$�����U�d��0�O#g��Ɂ1��@�D�&�{��p2
?� wx�l�H����W��e�-�ƀ�_"�+$k5�f�����:ӛj)��e���:ˡ�#8�����&4�>�M��� �Qut�{�K(��s�+���Pو;��?$=���\�(��*�$gQwԒ�g��4�[����㉧m ����)ֻԵѱ��@�O]N���(���(n����-����<`���o����I��E��������_�.�p�س=���� ����}��݈�!��Թ�>jqe���+-��E��w�!.[���易ٯ �/x����!�c�)"!�aR�k�Se��|Y��5/�ș�}X�ћ���Q��{��T#4���5��)W�q�M����� w���A�_�v˂?[cj�M_|�F��2�=Ҿg��0O�lL/�xS�s}D���Te}���ȟY�$k�
Ř����$�RHQ���Qz��4.�Y�`{�����}�iU��a����à�캝6��r�L�ʱ�ֻ���O�f�ɕ�S�:烃rܤ:!]��1u�������r���r_TxT$�J6m�kp�=E��*��3�i�_�� �2���Y�GH�� )b�{z�*E�s�H��u���o��}A���F����) ƴy�<���m{p�N�BQ���5��������XV%� q���e�J���_+-_�\:�(p4A��h��V^� �w�q�Ճˋ��ٙ%���TB��|7��J�M��spzX檚�4��uۖ�r�}���7����=�u1m>[�?M3�I�sOCY�E>��z���WX(Nb/%�žK�4l%�K�M1��$��j�!]W�O= b��!#��ry�3^Ǹ�dX贴�^���'��C� �h�F<��T�S�8�d8pJd�|����@���d��!����	5�ZK�U1�"�]�@������;�`v£��xF�+MZ)O�<l�)�� ��u�'#^���p�6�u�����"}�I�O�ղ<sY��S�4}���I����e}�э.)�I��W��Ͷ�1D��჌�ʲT/#3�����IC[0ݨ�Q=�����*�g~7=�ڔ*z0~�� �+�$��;u�1K��+��dN�Z47��ԍ{��Ga��ߟ��ZqgE��*�d����I���hFP�f��8���!I�
�Gm�/r{Y+���.T�lh\��h㈙�(���T��٧�M�K�����O����Q7a��z���l��u}慗��Nց��%o��(SH�|a2+�(����yݦr$+N��o ������]�B�s#�h�O;q�Z����m.gm21�D����N~��W�P�y���Q�UJJ�u�?G]9���ڃqK�� b��qCtL>"��9�d�2����5H���!2��KK�C�X�KR�	ʩ�d��F��<�me�G�%{�7=��T�b���gk��q��N���Q�]':ЁH�4���d�T�Qȟ��H��SvR�1W���S��E��ڋ5OCe���Y�[�R��Xjӯ'��a��Pe��=�d�K�X�m��2��0��X�p�L�-w$ē���3��������.��H�JD�?�ċv5�E�9�����*�'�jEW��( e�Ic��	%�j<���]ΰ�]������lPubB���ET�\OBp�n����z�u�7�q�Q�=B˚�?�ˬ�0)����?��WUj�'dȪ��)��O� ��\��n6!5ט�ވ��Ǫ�Xx�����܆x`�I�A���Z�j�n�����74�^�:2ֈJ�3
]��ro![���@ӑ�Ҳr�;f$�vhV|�����HHz� ��{�=�� �\�?!�G����1�-�́��w�8�����~�O��L�`X%=���ԡ��e@V6��Hۀ��Lm���F��"�B�4 ���%��%a"�4Sػ�S	�fa����X�mGɶ[46��p���M_�?�H��ڙg���P?�+�-�Ek���6,_w�	Gz{��$p8P���Zjfq%*����h��p����N��Ε�F��|�H�5�A�I�͜<��ᐍa팧8�9�r��.�0l�׭W���P'��I�wE�n��( %!�(�Z��6�^1Zz��0�� ���DW�g�V%��cx���q��?�NfӭNt�cE�����6�����*]��u�?��ϳ	nɒF"|�S�J��|��4�o����*���C5vk�ڶt^~��(4m���`5��c��0ad��f�qW6\��+����We�U�p*�Z���E܍R����,�Z�{ř%F������g���{��i�
��>>N�.r4���faJS�A�]�awz�z	Î�@�F$�_�2�^�(>�f�S���D����b�;�y��|��ZW�YK>��I�˭�"�jL�/V�QA��*z�t�+��n	dj�yt�yys��^u��
�14���r��3G�����ۧ��x���0���9�WB=�q��V����8�o��Yy���\,,���P�T�r�%�� \ׂwJ�bn}]qR�mC�>1|F;[�%�r���p	$� 59���J�%_���)���v�Z�!�Ƭ��!���ڭ���!�q��� >�P�(D�_y� l��I��`>������?��� ԏۓuǓ��Kj�����$�H&o|��K�R�u�e�Ԫ/2�fԻ{wy��TG�j��TR@��%&Y��~��3��x�7mh׸�P^;�Ѕ��f��@�υa�"weF�`q��KtE�G��e�F��/����{��� lbiT +pR���c�|B<
Đ�Զ��&���X��� j*�c�=�����w�Ak�3������u���5��ӗ����*�:�%�#/���?���{=_����	�{�ZY���ă�Z�O��[%�>�|C���ܺ68�T�FH�\+��C���\O��u������(;�s��H�#�d�E�
�g0hS��߶7�:�b!|�g��-��#�X$�Lt-���1�ު�Z[3N�3���,�k��(��A[H!lW��ѦEf!��B%&�-����4)K#BM���N�M�o�x��b��7%q�Z-����9��SxA$��yTz�������F�fP
����bR�a���\4�&P�E2hc��9F^��\������˹22'��+�p賽�����k'�ȎO�2&Q���:����4Xg21�YR������M��g�������$�mle�D7D��;:��=
����DR�xn��������=+�)��`<�; S��Po�]	�eȏ��6Pp�B�/�V��Nv*�
Xy3�K�4)#������3g��B��v�~���l�Ec�T-<)z)'��A�'�#e|�`�����p��4��<�:V� ��'pxY��UK5,!o�u+&�a���R���6-*�^�0T5�f��o'�Xd�u�{�Ԃ�>���pqLZ@��A���G[�8���T{�'�ȇ=�E1�h�P��b�����<^��ؔ)B�yE�(�0�X[�������8�9��`�[z�2��zo�OF���fuq>�?q���]Če��i�#�j����$_I�@O�^����Z�!�I�q����"��A�L�����V�Dމ�܏#`�[��+b:]c.G��πp����rW��7�_^f�PB�@Y:�2ٿ!��ٯ|�ŵ�����,.[ ���cB�/����(]%�G�M>���-�N�1��t1/�s�Ӗ�^��f�o�d��n�CR�(>KRĸ����Aș�:�a�p�w�ꚄETC��S�Gh���^;�ݡ+�R���U�����Pǃu��3ν�X�W/���w���˿�^D����Q~��[����$��f~�)��hQ��P�ԋ▹ʌ���4����L��k��,���n�'3lb�!(������mRm���o`#���U�P�S�y<��	�!��>���d��[�x
�NGv�����j�+6���ĥ'}U�i��oN�{%v���EU�8=;�����u�|]��xaBw�9_����!�/�V��X��6�6�
 �Z<r�(a̽wc�xn4gG����<���YI�4�l���s?{�#C��� ���J$�m �(����-�M��m����0'��?����0�҂�a��5�Z�\�~Ԓ�I���$���%�\/Iͮ>��r�L�a��N��nM�[�~K��
a��s��V�u�X���@`�pq#E1Z����Q
.�Mz��Tro��W�!+Z�;>�w�nӡ<��������V=���" '���'� <?$4ĉ�T�ZIe���J2Iq�S�P�`Y�⎌�w`�ҍ<���[���1�t�����R��E�}�A�&cX������D��v9R�@�fq���M:4(���H�j�QA�^Z}@Ga}9�1������f,ς�1OJ��x�EOb[��!$� B~I#X�MJ�&y�R'��>\Wu�X`�9��AOW��ڨ�S<\��j��t~���j#?�1���-�І	��w�L���\̎-��4���T�]�,U��MPg5�S!yJC�CI�X�q@��l<T>���a�Q#�P���߫��jQ�ٿ���f{�E���@Ӫ�g��5���ݙ޸t_ ��N�5謕����Q"UBB����oG��o���T�b�\����j�l���c�jnR��5jg��?G�**/6�ؽ��?��ۦ-w(�PP�LK���إ�8�7�*Hp+-��z��X�
�6����*�z���N|l�y�yT��PW���
�fK	r��:�+��H��,&�o�̧�C-r9Ac���j� V���"��01x��Fk�����s��T�[k�w:Acx0��a����YLm8q��'��A"�Z���Y�a��C?�*��<�۪����Ǘꆦ�E�&�r/���4c��$��@;���6�#���>�V�-�鄝���8Em�J#��F?�� �?��5�q�����|h�ԫm[��x���c�D!�z1p��4usQ�6�9O�T�7�� ;���� ����!7E9H��Xɂ�zL����I��F����Uc�?/�k��ƊYvz����e�� 2S�Wjbd�x�i�:�Q�J��,	����R�T���Ol>�rҋX�.�lu�{F��w�f�~Z�X+���-� Y��D�̈�sK�𣔹�3�z��RM�4%ŗ�5�.���X�J�c�G�h	�E���W��y1K��q�`��Ga��4�ybE�cA&�.{ڷ�1ߩ�[H#�Ҷ>[x��w�Q\[����������R���3\>?��S��g� n߃G��Ub���*ݝS B�¿c"���د��T4�|��D��J���mUa��Ρ<���Pؐlͥg��D���C6������X/�T#^h_�CB/���aQg�t �{�1����㐤6��yՐ�t�0<$E�����U˙Y�)з��Ȼ� \��OA��}���"�I�/%K�2��Ƕ2�Fڡ�� Ju����t81L�XN��5g�R�`�>T���k����ҟ8�Ѧ��/6�BF"4��eJ.&;��u�2n_.z~.s��#e��^�ߎj3�����C$��Uнl�_���T�`YVN�2u��V�+�J�vTw����;�;֐c�ժ9�c��y���3.m'u�G��WS�����3��0�ķ"��2"R�P(��C�9�����D�n�ަ>�2v��kg'���[�|��Cq���^	� ��YR�"�i��Z^�Ϩ��
T{M*z��C����+>��c���W�eT7�<�Ry��d`9�~�^���۷��=��	o�4���OMY�ΧjDH�1�
wz��	Sm�F/�j��r�M4�I�H-_�1E��!�5O�%:_�w.���ڍBS��]=��t��<���E�a�W5��4�y��j���+?������eK���+�R�������'�()�8|h����g!FU��[H�k�O�%I깳�Sgi�y���ҿ�qB���ڗ%<�[
�N�S��5��'��/?p������p����ygf�0쯚z����2�{/�O�	�=:��i���=#_,`�P�j���<c.X~�<|�~$�\y>\�������N��]�EC���c�g��Ε�͂�}�!Л������2$����'���6pfhew����н���9���ra���./�\^���VC�3u����#0~�&LcÞ��+�G���$�6!Ť�N�i�eZ$��R9q_��R��'��qʞ�ׇ �p��\:@p����x�Y�������Ż6|xы�U�=�8+O_,H8�܎d_"ʦzٹ)1���N�0�dj;BbK��e�YU9/�Z��Ρ�e��C	_�;�#�C��/���rE��w�1a��t��I��ޥ�q�ɉWC�8�UM ��K�lh�b�N%�r�cz4�=���u��������nND�U���ɋ�������F	���ź$},I�U���U,�#?�	Өzq�=��'1�>�T_aA�X����@$�5�@�P��t� 5]�8�ZΔ����B�jլ���9C�|6�����FUw��e����k�;��^W�P�˔�DQ��{Յ��K�5y������`��nx��dK*?`��P��XxO?����W�o^p�E�,�")��/C�����.ⳁ̙YĎ�x�u�s�����U���.H�]^-Q��ָ�mU}C*e�h�AU@dl3nu& x����c�����`]U����i8`�����o�-�ʘ�����iҠj?1�]��5c� ��zftDg��_*�!��E5�E��fP��e���7�w���+�@ïZ)�> :Y�VuuC��� ��{���,&q�y����:>���@�uBd�(�)��BkA!��'��]J�/`���9c�B�R�(�<�Y����z��(��.o_1�z�v�6�]i��P�ITQgյٔ���D��i#�3Q�|�ZN��n���'h+U��������v$7N,((�(����M�c��m�5����P����֏.NO����k�o����ң,rm�J3N@��Hl��OŹ2��:�]~���[�?����+/�ƽ`̚�]���iD6�8���G��c`x������z��x�hMbœ�i�$6E��x������'axrL��~�V:��-烲N��3r��}�)���8�ߊ�������l�ğ�}�X@@
	*p��#Gb�T΋-��;
VK٧E�3�f-��`)2�uX�ͥ��0~����$bb�+*c�&u��VaM�ow�K�������'��vϐ��GO'���s�|2��l����5�lٶށ�[?�J�c!v�{0'�t�:������U4�3Қ[K���H��
�� .߼��Zu�zHV�t��Jv ��%�|98�͆=��-�ާ}��:Q=a��t��C�O�L}�A�a�}�7�4����k�9�l1���aM����]�5��)���F�V��՛,D�]� �f[���͓A���Vܒ��`ۙ0 m�-c��P0����֟5p�g������a�*	τ�D ?
���ed���;��|��zϬ��c����?��(���i{����{n�jh�v�n2AƬ���Mx7$���z.A9x:0�����f�;6�#�W�*Ut��F3�����">��Iد�I�Lr��`/�M�����G��%/�ҋ�_
Y��p�,@;�ٿG�%��]�,��F���f�7o�.Kr��"�'����|`�OmV0�p_�򙚅�5�xA+Ζi���8]nIb�d��̜�(KU���+f�����)�vvZ���)^�)S�{�e���Pp�K�!t;g��է��p/ �:~��j�,��8�����j��m����	���wc+00�>f�����wOێ���==�r�'ɢCV��s�XMJ�l��צj�粷��*]�u����^rDa�{s��䅋����|z�{�%$��_�$��)v2�GS:ؒ�#}�'cbT_l�;�τMO������}Y� <�3�6���QX�ѡ!: E�y,��G�AQZP���Gt�E�6��w,�RbZ�%��/6�L������_[�j�D�	�X�A� ��A��P�L�[����a/Z��il�N~J�O�yZW��jy�װL���m���$C��(�FN���p�{�T�A�
BM�`=��	0o&V�w��sr.@,�@k��Â7���������*b���t�O����� �)��n��*k|kux޾��Z�T?���y|�$��!�����Wz��eUO��|���U�3�k˓����0�kK�%ũ0��=�G�U�	�Q�!�/y�e"v[�l֗�۠�=�.�)���N�P���t>M����T�3|����2�U�9�0������o9z�lh�Bj��`K�]�N��dM'�n�_S����[w���98&W�^����cgi$��}��eZ��Pd�5�w�ۚ�]���!�c�L�d�,�S��c�GPK|�����ҡ��e2�/�)��.�y��d�w�*Md�Uqb����W��2Ac�z�_W� ���֧9&k����M��&��H�����Ť�E��`�?�΋m����ـ@:#�I��̿Ǆܥ�Ƚ^������`�nE/9��+I>�\�x�1._���+�أ��9M���{�r��V�S�K�^��`�A �}��d�F�|��X�+^���:#��p&h`�f�\�+!�>ҏyʧ�3������E��9lV���~���%!?&-���� �vAh�m�Řy�P�u��p�lk�53k��v9=C\{��f}��`���Z���6�x~I�Z�XH�.H���b����MM:����M�Dj/{y��]�^���������fQ�]^BL�)�C��[����m��E'���Β�L���wȾ�T?��qa����U�~�?pA�R�Ŀv�곩�An�G!��i�ټZ(��OW����Z�)r��%�%T�	w�H�U�ZYn�<H��/j�kn�/ӆ��Z|���sPƊ��ƔpL�,����ߐ�1�. ���q/Y�kd�7�ʻ�uҘ3�P�
�J�T����]޹[�U[�������ی�K�2_ k@H}m%��,�Ÿ�ܨ�^NF�Y���rB����Q����d�?&):�ZQV�tͧ��a@���@^�i��%Cm�\�)����cgY
5���Y(/�Ul��^�5QǾ���縴�4�����w�H��O[���%��^ �G��꛻6����y��Q���L�������;�už��*�u�j�D]o�B9z���/�?�[t�@�ʁȅ�6	��2b��O� >��p�* ��:����/�|�m���Pgu���v�q0�)��ې�$K9�����?�G"����"�aӢ���ɥ�'�-�c�\ aK$��bg�ɇW�ń���ؓsM�k�I������fJN0�����"��D8�m�	`���I�R�����K�8����t2Y�c�/�]K\n��)7�6(h�\!c����3�H/f�y��	�ؐ�݃#����}J\��au�nL[*���ĩ=�S�e�~/#�Qi!��C{����m��V� ifpE,���ϐ�hԏ�^?�N��-.<*�[�c�%�;��c�����T"�Ñ�%:φ��	r$��e�Gpn8��m���N�{�!�(J�@����3�rb�R=�)�qE_��ր!r�\�c�bE�����>!�G$ ������q�;7�(T�0-��\��&6�9DFS��jr�k�m����j�t�-��P9�,����+���⽶�� �s�.�.�8����UO��C����� ]7Ӗo}��y��j{�6��6(�[���n{b�OHC�C��{�:�E+����$��m�;j��V_��r�<���'�؄�xHgj�ބꐳ��붑�Jv.����������c8LH!�
�Ibr��Js�ۂR����[ %h��uH�f�e�Q��$,�:�ߜ��-��n�A�0��mM6��� 	�A�q.���S�5:f�܋�<o���vA�3ZT�g+�W�ς�*rtÒz7h������]9~�Ҷ]�z�1����]�`�-�)��	:,h�n�Å���VTxJ+0QO#�X)�xN�R�"Hx�������B�'�\�V�X�v����$�?Nb�Cw2�k�.�����2�%�t�Dӹb�~)��)��y�Q�����0	�\K�>Ģ-�	J�gY$(��R�m���(dPNI��ެ&_&,���.����˺��<ݴ\��A�vW��ӵmb<q�h���I�̽� 3PNW����4b�T�ǋ+x�G�@v�6�uhɱ�~�KP3S�H`��@��V�Q#���^�L�a�3ț�(H���zǈ�`jS�]*'�@�/]�40��K��X���_0�Oƞ��"��-�s11�0���n�HZ�\% ���P�R��eق�0�v��s-W��
����z�������I��G*�#�Y�������oiB�!a�(Ӊ���i�q�ctOC�`	
�AY$*G����r�="X�Il��PHҗ��A�N|�� �42��p���j˶��\��n�{(�-|�g�*2
��t$h���(�}��^Û%{��Ȫ��v2# ��:^V�%.�
��5������Pu�p������3�c%R8RvkкGX��d{M1/g��7�X4����!�nU�c� �^
����[�P��,�kS^�����]R)(�tN8ȗ^օ��T�"n[�p���W'��}#���85�H�̷�璿��1S(�i+Vg� ��8nq%�_���5��k�M���0;"MAbd<��Q�(�����{�a�\}�[��ni�F�����c&g�엯#���Z>.W��ߗU*e�
�%�Qg`�|�0vG�rYC�Q����{�g�v�)%��_O�
,"����`N�L@��4��\n���,��5BM�o���1řea��k��XmMg�_/���ժ��������ݓD��ߩ�dǃ�����6K�D(X���Fcl�f�=���;:���L;q8�	a�}��栟�A��:ʿp����_X�Y����j}����%�'�� ���a�TD������SF�i;o�=hy��Sxk�O�������G�,Kmlo���������ʱ�_�Ih%����ͫ0�a�ۤTW@��j��AcX��ŏ-��.�-�:cX�KE��n����g-}�³<�-L��u%J�P8��x�-�=C���Y� �_�R�^����T�U��W2[��U�cֹ����n�.����^��ŭK̜�鸚�r�4H�N�>j�!��f�U��nؽ�K��R�F߬�������i�Ш5�����9�η�/[� �o\��ANZh��Qh1Z�(x_BS��{]-�Z�b���_]y��M'A�M)/;�oO-m�:9,+���4�ʅ��+e�d���s]�6��T@�@<h�/+>	�F=x�$�u�p����3��%�y!o�����9Xo�HƟ��g#��.1�$�PRX�n�u)��[���l=@�C��9�������|� �`�����GqGV]�&1���"�衖΋o�1?Hkԕ�x6�D`��|�?�D��zk��MϚ�Ez0=��M����2��є�,踐۔Xg�k"q�[��7~�N�G򲐤K=�A�FZ�,Q�=kV;ӳ�!ߌs���q�p\j���80�1����M�Y.�����S��f�z����m���M��+D��6�I;s�`���0��������p�t~��JB�:=ՍQ�����`
J�Ѵ2#V�:s�F�b'⪄�g����7�0���A�w693O�1���p����nҏ�G�����x% b�4v����e�� �2af�:*
��������h4Ѷ��������sL��Ĥ/+����`�r�7*0��v�ť�h��
ĩ!���<x���%����ilU��J�}�W��F�m!"dƣ@�K�	f��ZiDm����f�4�+�s��?/g����~[�P�$����	T�١PMw����R���?�,����z��o�f�V��kH�	���R���<R�ꓗi�#`V�v<������-�<$���R��L
�c�w�Qi��\�u��B���Ѱ�4N�K�F3�rC������e���@��x�s )
��چ/�9Hj\=g�a�I�@��b���F�ndYDb��C�>d�����wn��v˛h�j243tt�+]���B��(�E~9�I���W����R�Y7���h� Ԩ�+��[��1������g�<c�1�q����8MM�3�q�ŀD�%^��M}��,��$,��r!���vo`�`jG����&�ٹ|����kn	d'b<."՝�{+A������Ha��뿡��-�G�����"��@.���CSi(d��KM+�]����/���h�¡]�P׮쌎� ^/]�"��C��34�B��:���&��>h�gj̢L�r�Y�J�t�E��Ce�u
P�F�_��j����o,�����\�}��Sa�[#�%A�`C�|����Ïd��^{֔;+U~��e���96��o ��'���,�`؈�Z�V���@�l�c��FB�J��Xt�qb���
�h�Н8��w�B��������W30�.iUl�)���߰�HX�Qwt�Ǒ�b�!.+
!O|{U�H��RY���#7��a=]�{��.�=y��R ��]�zm�f7I�m���������>�fN-PV���1�S�.�ȝ�r66ި�"��swƯ��'V�C��P�Ȥ~���1ц�POՠ�~��n����.�o��:���0*�d�ENXS�5[�R��� W�zyW�~�L�s7�	E�4�\Ij��h·\L�=�4�gXEk[�D�����Tu��a
q�#~ZiGK㑫�֙��Z�Z+&��ә�?��|��4#t�pqA\��^5>g�� ��$���X��c�n)2p!�O⸷�'%~�RH���g�l��R1��u�6��3|M�g\/�gT>��O����[��^��L�b�/�;�� ub� ������P���e��,��K �y=�w�`��������v���l�b�~�!W,t�Z4�2!��]BD��9brH�o�����4Ϥ�K&[?`�Tb����i*�)�v��q�bH�ϟ!�tV/�hd7�i�ç��PWE������׸V��F`D�I��?���2;���|�� w�Y=Q���3F(��r,_N�%ݡ#x�lqs�<n�N�E����=)��j���zVYy}��5���	�襖jCs��S����+���do�;�_Mc���� �a^FM!v��4�&�p]�,/���J�� "��;�,ht t��[�۩PP�<x\3A�.=N��&)�� х�A��e/"��%���;�� �����$a��YÆ)��+�X���b�}%
�h0E����)�E��:����å�G*(h���b�ֵ���~.K�yE/�P���KY=8u�d����{��0_m�r3���Ϭ��,�0���wT��B�������@L'�:~3���O���7��!^Y���IoM�3�ͫ�&!�E�������k:BN��lg�z�`]۩Bzk�	��o��7��jO��[���\�ᰤ�;$u;/'�b�B~H�{C�r~X�Ƽy-(=���4����]�SɄ8s��U�1?]�×(�>��m�L�&
 Ӹ��y�y�mc����u
�n;�iۗ&�>���"�Bځ+�Q����e���a����!Vpi\֊W�'.X�S�>O����R�t�f"��n�<��q~�؄ئ�e���/|�=M@V?2��2�����ž���RA����@
Af�`�Nbox<Z`�mE���}�{�ɚ��E���=��P8 ͟�- z-��o�J��蘠�L�!!�A��_��|�pؤ����ՏN���-qS�ki/N���ҳ�M'�`2z�P�f��ԗ��it�}��FE�i�3D'b=з#?lr>��d����J����"\�W@����mQ��M#V��K�4K 8cx�0�kn���X7Y.4�P����u�N��8򂪀6_���I8?]F}At�F���r���+&�q�G��0V�wAvӂ�2�+Gd���L?���z����o�Ѽ���`�;(�q,ȫ�}ٻ?�;k�@S�(9��^ǳC��5?��{��V���%Z���^���h�rR\\Ű�UQ�s\F<q4$�lp\˕��̘���ɝar��v~��=P�ٱ^�8� c$vaQu�S����gJ7�z��{��D�;�|����Ǚ��=@�Q�8���$ZϤ_����`*RO~lOK��Xr�;�y��(�Z:�����d���מ�/W�h<��n�4���y�k��X���
�B��C�1j@c�;�����j/ݴ\�tC>\%,M�Sg�}�U{�� .q�Cy�F-�Y%�	t�Y�v��j��d�.V���M+�t��Y�?Ĵ�w�9��n�p���c��X���Hlw�+ϵemG��<^�����CV��{�K��p�x&�'/+(N��B��Tl@~_^�{ʠ_��ߚ��A���J�g���yTs�dmma+��@��K�WaQ�I�q��<-��ϡ����wy	��"��ΡώPB��?� �m��)��?!;'A������Iқ�,C��;�����6=8d{�����=�{,e" 3��x>�\��NfJW�J0���*wQG�&�������h���
�91���?�ڮOK�� ���.;�%~%}?c�V:R��P�!�������)������W5n��[�ҁlCSZstb,��qM)6$~�V�4{`������4�gȵ�q�6 �,Tl>
��ܰ-`^Q�D�GN��Ü=GF-�C�>^3h׶:nh�jD�!7mi!
GƳ�*���t*�\���])Є���sr�I��)
���(��C2n4�_���|�-�.�A��(�l�0�_��%�g 2�n�*�\D���e��Z@$;4��`6
�;�}�Ew\dYg�D�;�N =u�^''��y����&T��#�� �H�7*�7�afY�qH��t���QKsiMՂm�@d�@�J�9 zK.w���G�?YA�q͕͑��C�<ʋes8�#ɽ[��!�+ؼ~���b�%���*�*Zg���Z�	t-Eڝ;��!��N�Z�l��~�k�h���y�F����)+����q��lV1�F�B�>��mP��H*����s����%��Q�O6��&�cFg*z�ڴ�Ւ�Y$�i���;�P��._�n�JB����eZ�-Jw��&��_��-�JF��"�;�@�j�4�o���,K�h���]����jjl�m/=�;�$TA�$Pv�K����n6��;O�۪��?��zjXH_ɴ#w��~��]V��Nф����BUD7����S�� F3�P�u �}#ζW)����@�}�/3���\E���2^��:�C��M�����bbIJnC��%����a?�$�RGX~�8q�mr8��ך�h����[� �r�F��*�y�
�Ã�8�**�{BC�(DmWg�t�N�0�����G���u:���z���a�_H�W �(�Y?�&2��QZM'�G� �0u���A~���NJ�9������f�m�S�M���י]�#k�׋�\xn����C�2�e�#kt�ݿD+��0S�Go�/g���}u���5�[�L�W�<�;��W��{e��ܜ
"�n���=�Q��a��H�L{�;�X���!���D�UN�R�l�{WfZ�� 0�N�Z��ǇM�f�4�7b�p��_e��*껖����|6A��3�Ėt�R��Z��,�����0,!vQ�(9!����ڡ��$!(��u�o���Dk)�Eq=�=n����n�4��['��hl)�
Ys�.�b���B֊X����+�\�YN���r�M�@2W���������,cW"_�69�xb�UVr2rݤ�;��}�׿]@W#%���F��XZH鬛���'�8�֫kǯ�˽2�Y�6�ʨ�<���vJ��|���%�cg�4��Y�{S��������͚���T��)^D�ܙ7u �rҺ�[y����Sw�S!s����M��ᕼ���.8�N!�1�a��<4ս51��Pz�<�q|1�m���顓o	��1�F[+�w�1=efӖ1�B< ����Ÿ��H��?FN$|f������i.��p�8R�ߐ+)��	N(�f=<6B��n��e��R)��2�Gb�C����1	�j}�a3�ga[���ݩOSî�:-��,ZJ�:/H�^g�t��H�/����7���J�\�Z�͈��?v2��Ъ��+h���I �D���4��5��x;����\C��]|��!%hZ�t�~�ĉ]-�\��j�/�խ�"vd�D9�^�Z���̮W�X)s�X5���D�A���TU<�o���6(�j{�쑜BP%%T~�Ҹ�p���w��^�W&P̶�hHr�e��b�z����.��ܛpаP�u�}��7jֱ �����_���6���Q�@��/�/:��1#��3�#���p:!�"Y 9b�J����D<4��2��{�d��bR$��֖V�I �ʬ�o�Y�pL��Sj)^k�K��9=ǖ�g |LF�2ݴ=�.�U27�N(��C���:�aa���!pl4��̊��+���b7�[�K���x~�l+��CxBP�������L	�u^uz׶��V��u�3��c����Bm�WJ��P��:[���[�m̾<�\?Կ*���|W4�V�${���[�S�E�M��Hh�4��/^�y�d�T�ݚ>}��l�2
��u*Q&�����6��4��TIVr��ͭMD�����܉6����>'�U�����Yƫn	���H"e��!��%���(ޅN�N��ST`�{m]�����Q���ƈ�ٿL�~b�A�z�m����|JA����W9�I��)��:���z�ƬźF_T3�� I��ۼ�
�����_ng�N��h��OVc_6��
,\�P���P2���㵾犬����4��Pc8=��c4>Ð���P�)~s���4[ʟ ����Ś������Gm�紼6 ��,��@����\c$5����Ð���b�4��%��I��"68s��@ ������̳�B!u�2����*^b;e�Ȧ�K�٭l�O����9����#T�^�j��Ϲx��n8�l�ƒU�`DA����h��g�[�Θ 8�NF�\(P"��,Q����[r�΋� ��#ƔbX���3�4�k�m��FO��K�����!����wjE�-�e��]d��{�@� >��6�"���be�r�����1��)t< �� so:E�A:HA[|I�i�DðD�w�K3Ѹɭ�|,��	%t���p���9�fj(^$�U mA��/��ġĽ��Č[��A.�D�Œ?EQ��/n�
���͟񄙠��)GW�����:4eY�	��v4p�O'ѪWH{F����V���'|��z���Tュ�=�pM�C��r�ׁ�|c&��#V�>3:����J��
>n�D�Gio��8\�.i|\�Y �s�%��@AG���}���R�Z�~�kJ�隲�9s%��+���iG�u&�ލ(� �>�zv�K���C;��3��r�o���s�&-Y!�F���㷭�̗ЃR	�e��؄��a��},6G��b��P�:��	' /dq�C��H����6ʁ!HZ����<#̅|vk�4U��ivE�g�]@`P�6��HX~E�SΎ5�xS]���9�����I�)��*���ƕ�SoL��8`;W���O�ɐ	������~0x��&]y��l��l�c��NAR�s��D�w�w(� �3��JO?D̬�Qσ	�?=�B�����}N�.U"MT��<��0K�K��7I\�}�a��:���ۖ���PUE$��%R!Î���n��G�_p��o� �ԛ����U��P�}��\Ƙ|@�3T\_{u�a���T��?��\�ڀ�6[/��h z���p�<��/���M�.l�*�N���2h����Y� *�1���C-Wt���y���N��/�&�v܄ h�jI�2JB�j� ٞ�7	�|��#	,��Z��q�(p֍�ql����
�q�M~��+D ����R����&1�7�ثv���NV��7� g���N���s��_<k�%u]#qrf)V�<��e��:�P�kL{-�D����Ĺ�=�#`f�%׶b��q� ��_�v0���_�W���ċ��9��-&,ku��l	� K�'I��������W����E;�KX���ZҜ�#�6ÿ���ɭJ2�2Î�
�v�L���qR��;,�:#���k�mH�, dF8w'z���feݮRM���}k��_X]�F<���x2qn]���З�8d���i���%�k�9�2�qP++[.-�z: q�l�NK2���N6�x[�>�ؖ�����z��`1����8��ۂA��e�H�76y�~;*CF�Se����p9z��D��]{P�f-դ�U ch��E���cn���
F ���;�Ē�}r=g7�:������Ra5���~Yc���_W�=>_�]���Vk@����L�%�WCo�E��>��B9�u�������sގ��-��67��0/�'s��c��NPg��d�83�āiū,��j��GnƦ����d�HK����q��X5+�q���W�D�������=4�<��%4c��c;[�x�U8X,(�/!kϼ��?��;j��wFb�$L�^D�=�1�R ���	Ws5�d��cm1�5����R-{���<�TU|����sΡ����ݱ:��a�T�����T���l	ܤ�{Y+)g3��%_��PO��u���n�-b�4T *���.?y����5�1\P��1�Qx���Yoo���\
%�<���IL���N,I%��u�'@:�rg�)�iǬ�����N�e6X8��oP����tzc�� c|Y�6��	��̷�Ֆ������a�Hy��k���Nř��8�ҘK٭�O��%10��$+{^;]�i�S���$ee|��vsF��l��"9����Y��;:�s�+G*�˥�T~(����MZ�S�[�,c\��R�n!a�/�3��g���BU�!��h/��#�)^1�"}�Y��H��83A?��w��M�|}Uzv�X�p���PG\�l*������p2�tJ[�x��;�_Ҝ�s�v����s�^ɞ�����nL�!������.�KV���kw���u8)�j>J�����kY�h�>z*u,%�r�ݟ��\��j>뉆^W���u�j�sT5t-�)�k�O���:�b�mh&K{M͵����6�����N:�Y_Ud��*۹�Ҡ�y���=��n����J�y�<a��������v�$B��Z?�`&����28�<{$��93����$dF����?Æ����3Մ�GiY��#����M���fۀ�L6�� ��jd�Y���.t����MY�V(���϶��ZAvh�#�`��'F���sT")3A	�?Y��
�mL7�^� ���Q R�� @u��I���a4+�ĩ��v}��j�J�����e?W(���c/8�X̫�۾��~����)�v�"����塼�\��9[u�+b����K�R�6_���oO�U��$26����_:q�:L����H�$���&r3}���)�z��k<��Ƹ���3L�?�aO)K�0�k,��:~%1��̿=�ܶU���Tf_7�| ��t}�j��S̬\�O\�JX�p�h�*���_�6ɿ�r�:b廯@j�v�h�z�0=�9��-v{���7��^>��L�����~QfU��t�Kzw��I���o�z���ti��h1ՌjFT�{�5��{ն/Ez`fl<~M�#�nő�W�fX�Iq&�_���B0��3�8���xl �W�RJ��[ʜY����_�Y�N�X�:�h䗹�"mR��+�;e�ĆsPx-�W"�}gt-�rG��*~q��n]G��J:�5���gL�D��W�R��mA-�֙��ˉ��k���MH ��:���K��=��Dמ?�Y�����x�&��3�4��ġ��J�6�X�h���t-��p�J��MLy�y�vk�S���F
�B$ߗǬ�4��3&Ғ��*�OпF�.��W��r�'K����bx��_[� 3��C5�����J���{�se��(�F��0G�y���Ⱥ�ↁ�t���ڟ�N��orASnm�y������۫�5<�e��~���)[��]�SzY3������+�aE�6
��]y"�Ѥ,z!���->�s'�'���[S$�u[��B�Y1R>�X��f���0�%w�RF2��aew2�}J]��Rv?�[�O�>��K.ª ��3[�c	?������ȅ�<d�й�/#�7�@vW)Ek��nr v������nDJG�kYy�x�(�]h�wA�瑂��%ݹ9�"�O�vۭB�z��#�G������5� �5�g���g�&=�.�����|�N�k4��a��{�0\���䚍��H�;s�T`�]�c 1^�
��L1�\S��Y�u�,�kg�!�V��V��C �k;n[ي[q�6TR!�B����KY���?�L��߲��MZ�y��py�V%�-�DY�%w�E�k��eF�R~� @�����ȕ�Y��6��)tWE�T." �@ u�-��$u]�B�	P �'�"��di���oo_Hɢ^z�o����v4� wpNM��5��I'�P�	ٞ1�����:esq���h.�����\^�,r��y���JB
�jY	��U�(Z�w���Ӣ�vlI��o�9fd�ϭ�{~��	k��2SE`��_�d%ȜI���6oU�{�Wp
��-~�<=*��1�b�2��2/��������$<f�i9��(�j0�~�V��Z{ӆ�M! ?�v7;R�J6�7�%�T;G��<�f��#DĹ$^=� �	[�$�Y�.�? M�ʷ�GX*��3p@�	�L�z��u���c)�y�xb[���;(V�@�/�*Zul ��i�p'R��7����D�i	ʐ�-Ū��=���&K�V4�r�*;��Ń�A���_a��Z1j�ӿ8w�K��L�K�������ӡi.�Lp�i}L����EuM���8}��Th�Nȴ���[��N�n��<�m8%]o���FC4Hy3�%��F,jЛ�8D����y��l�/������#QY@�5������a�3�Z�&�V��=�5� �Hܯ�$Cǲ1I���,�Uk�� �;~o ��R*L��@��9���Þ"��-�/L�9���N�c7d��2�#����V�
��bwSU�8�`@���H`���4'D�Z����$�l�������g�#ax��11�c��qۦ I\o���c����{�`;��UאJ.������eqYd�Ů?:��h���P�� �(RISF����ٮ��Yy�{��X�ȼ�V�a�Qs$�T��Y�h�})�+]��,��UJ�����&"HY�e����Ξ|=�h�����u{T�y���(0h&;{:�v���L��}���J�k&���P�Ns�vox�-��ϖY�G��{B�f��g��=B0Rj�-�2�_�L���XD2դ(M)n��Q�(}��t�PD�L*H�J7�OUrY8����2����"����4�J�п�ucc��6�H���7̓�C��\������3��$3$�cka������>�/2].�����,wO�B�� Y���n�b�R�mʾga�Rpr INlΤl��K�%&ȭ��o%�Uh����;mVX�`�wmt{y|�]�,��@D����`���9�<�����0����Y�9�bAT�f2R	��4�-Ά'q�x_Jue�����r�@6*�?��3-%����+�#�r��Y l�GY'G��07	��o_��=��ͅ�P8��Lk��u|����pG�t�p_;�%���X����	mn�!&>X05�!��Y	������.�����:q�"	�8���_m؍�4M ]�=����]<�6��R��{g"(]2�zʳ�R=�n�B
�Ԋ�Y��ȰT
v����}o�#���>��#�]pF�1c�7���V�dk{
cF���?ä���Ee�M�.Ͼ��i.;r5���B���O���'=�_�����,1=�01W�r���(`���X����ʑ�ThbF�Yru�G�q7����jذxB0�x�M�R�l�~��*ك��{�ό�gF���l�ˡ�U�¦�K�A������P ř��._GWO��9�ò�ۧ��oP8���ubT�w�7��6#+��{Ұl]ybxQ쇉T��aU�k�'z#?�%jL?:�Q�h�O�����!�4���ڧ����BAѱ	-]-�e�"���?��a[�8W����`{��ٓ��廹@Q�ɜ�ҝE� �$V@#���2}�s��������)��H�~`
JTP���c s�C�-W0�Q���&��Tn���呼"ġ^�:q�	�%�$Ug���UV�G��i�LŷR޸��,�a,'m`h�˄{���4�v7�9�-�k"EX��N�;���y���J.�A.� �ܖY��Qpub0 �4 ����\���Jt�[�ܓ+��=w����GGD�UY��Kq�����{��Y�C��Cۂ?y��<��p��L�E!��o>��z��4��z�5<~�����d뭣猃c�),y���E�v�٤Qe˓��5?��������)i޲7�/`tJi}�S�������ɸt�t��*���JQ��Y$j��x_}i|2_Y���d �����9ӕ��K�W��(�ɳ�U``k��rϵ���Id�_f��z���?ְR����d]m-K�2�i�:���@Ǌ���W��/�X����9����6hB2FV���L��?o4D��jW��5k���N`�C�4;���<��<��~D�3,�8jl<��v@�"wO*�[����}�|3�&�J�ɔ�6W.+01���G0s� !dB��	!Ar�M�=�Z�"G������e���܈z�7��"��b�>I����`�*&��`xS���p��&.��Dyg�Ы��ǖ�%A><���oȞ����Px�\�k������,S��*�v��
��;j�k�b'�Xeۄ�����R5�QC�)r���%����2rx�E�R&�CΘc;�����p����rD��<�lvҿS�s ��M��4���aą�Y-�@���mp=���8$�ǰ6P�穟U����j�j�����^�N����9!6��nڪ��;Cx
�T���phQ~a�b�D�˓��g��>�$�<���Kv�\�cO�>��^��B[Q��V�b���pu�!�zɲ%$��:�)B�F�z�����G�r�]	R�y���7on�&-b�1��!!����4�n�T 7DD��	�'K_R���O�d44aHe�ȂvH����d�Z����7\O��&�la�!Ɔ�����}��P� �J����&.��s)hav�J&0�!��I�y�fn�l��F`*0Z�uj'v��ʬ8��������r�):q��{�����v6Sqܕl���#"�ۣrGt�KO<����m��q�I��0t��x�}`��7f��sGi�u>Jѥ��L	윸�=Ƅη�?'M5�3QH�}ȿ^lh���}���x\�-LmD��Q@�ԍ>R��4�|�qU�ڞ��&��k��^ O�Pĩ�P������i��>��'���wya�(�]t7�pB�
���?�JHH:gZ彻N���ĭ/oe��fͧpA+ޤ.�?]����i;���	z���l�k���xQ$g��oH��<�������qH�H1�B����b��=O�#*��L[�G�RKx�~sm
�����Y<������1]ۆ��`\/G���7�g�f6�kyav@���t�$���>�����X�PEX1�g"E7�	�U��Ny�l}��=��뀊nn�߀��?��P��En_�c�b;S�fW�qWi@gr��#[��}��N�sh�:[�I�tk�L�RD�1Gd}��eSܸ���?[JMӭ�k�z��P�C�a�N���2�~��7 Y�g}� �^riT��;��V՝߀N��唫+R����ӊ�G��7�AQ�	զ�;�C;T��!�h~�F�<Q*��ş���P�FaD�{"c�`�]�4ݎ2�US�ݓ����Eɬ�jc���{��а2�z�H(�v����1��J%؍�3
��y��qC��#;�2�O�PX#����H���x���0��a3'Y�Z�H�BNq��Y�B��(@�� ���$囂� H��C��<Yv��\Oj�I�����>���SU�H>��P��w`QuJ,�����O�Mƅ�?ͥ�<co��:A�h��0����?���S,p���Al!��8ӷ~�)	���!��X�O�E��$v��\&B�(nF�/5��KLv�5�3�"��:e:K����`����z�!�V�������(�rNt�Y��'+��1���V�} 8��TE�s�#�
��=v� �Q�R%�.���a�L�څAV�i���u�J�d�Ĥ�,���`��DI74�H/�>���4��䜖�|�Ѐwd�g �I`|��.k��x� ,����� ��|���p=#��i�j��'�[B3��3����QO��nyz�J4�W7��W弞5�£�1�/������q�s��n�X� �Bз1Gض�B;��~�9/A��C�Y�\�謊��I�mP#�׳6�;�y]��K(z�j�?�eBR�ů�g�3V��V��ZXlgъQD��S��y]z���
ISPHuG?�>Pޟ}6�%����k���69���ԥ��c������W����ϻ5���?�O$�Q����='l���X/-��s�#E� �[۲�a�P`)<lqV���B��	��@�"�0<��z��|hhd��ܯ��Dƪ-�;�e��t�'��G��eb/�˚�g�bЫ%� �m<�����F/���z`���<�#c�yN�c�� sߓq<�ԦC�[���M�bqw~��%g-)�)�U��+��j����p��6��D?�ROMLm���eĎz�*/_�&j���B�x���Ù��=��>fz�o�8�
�,���	V���m̭c'��)D;�a������k
H�=����&�}�Q�*<}�{]YУ�i�Y�t�ʚ�&t
�]h)�F�G��a��m<MW�y,,��[r�I/�,�Z��ckӲ���t� #[`R���1��m����9z�#�⒉�s�����ge&=ʠm�����o�,���:4b�m<走aH�{���6J|�9�9qI���ntz�UN�n��� 3�R!$W�	S�G��-� �"��-Rؖ>r��~e|ݡ�t�֦"���o�7��t_̼+��=#���@2�-�����;x�/�x/7���Tē�B��kL����-s�g�M�ԏ��`l�#�y���a�>� �
�hM�ճ�N5�˦���E{�z��ω�@W#�U�vח�v��U�d��h���͈{P;e��ͧ��~/?�f��8��l��j�ϝ��F���{"���IPH�t �m��?��%w���੶r��OT
������W� �R�d�j���ge��ZO���40��-�{�#�opSg��a��h���@W��%���[��,2Vʎ���'#��C���Y�Z��	$�V,浱@j�㧜͸+�P�� Mw12�u�������D媹�Z������l�x�)l;���0\51J^�gX����[� "�n��=m�#u������ȴ������]���!�VX �=�x��\�{L�"[��S��Ci~)7�����������tǤҔ	�?�5m�$0'̹U}_[���0F-w����GVQAmo
����_��<,#֛�|�1e@�6/3%�W$Y79P}���0�x��Yc�8{�o���$Z�7��>�T��+�_�E�H��VH�u�B�J��<����%������'"\*Y5����O_�Z�60�(�y��3X�ic�Vh[.�a���\��$�˅$���D�?K|�>�$� dT߁h�-f ʻb�91Ȫ3xl���D�.B��4�Z|!SЇ4��+r�6ll���
6��6�ehgEye��U��s��%�	.8C�,-�Ҏ���]�n���?甊 D���A1��&1wB����=Ixd�0��D����rO-s]C7V��E��[ڢ�n'1�i�4\�����z�w[e?K>��N�2-��7�'"�D�#���U�~!�cV|)}�]����U0>*������r�T�'���8Lo����<ck���:a��܇�9�Llg�4�$%�8�E54�y�� �=�j�֚�-���d�ǌ=,���86��@�-;E�?�w�ĉ�Sc<W�y.΃��n\��RMvТ㵉�ц>��E8��?�S��Z���?J]�����?��������U.dYgn%|�a�sq1s�&i�\ԺZ]tIPכ�%�?��XN�]`7�I.��X��#�[�t��b�EJӲ!�N:�7>��y*�����AlW?q!_�M�h�w�A��~*5;���R���u�g���Y�s�mԟ-�/�K�><�"�� �w&�g�8\���s#�Z볐">�ՙ�?#y;��/�W�a.�~�s[�34Q
v\�+$���z�q� ��1iqW����*d���z�@ I�
�W��~O60����f����࡝x��xm���0"ʶÕ��8����s�=S#$C�N�Kfe�x|�ٻ�oC�HK<y!��xU�x��y��������r�Ҥk�;����9]y-q�(ADHT1(p�
��H�3$DW�;Ѓ{�jeJ����%doY~v��ᄞmLJ�jk�Lc���n]����6te�@6���ל�%�H+���W��>D����B�;�ǒ�o�f^hp�֯92۔A�ˁpN��Vpo�<�}k�زu���(y�V��b<��7�X  �<'�Z2�A�~ F�O��*���A��RQ��=�E��;�Q�wG�BK���aa��8��P�^ٞ�X�b���NӞ��q�b6W��s�M�I�T����쉧.��ΥEC��FI���)�P����7�5�)���J�Ev�*Y ���h��	��'�͛u�p^aS$���F��<��R�(ڤ�2���C�\�&�6nm�]X�Uv{Q»�i^9C �4���p��^��O�q�z��+���XT�� $��$��.�pfD��&d�~��^/&�O�\����H�'\��'�k�}-Is� ���[���Q�%��n��!�A�1�a���Z]��+1�����yJ�al�F����9�\�	�~l�;���)�L�����,�] ��&ALq�E%��Xq��7�g�ȁ9H��u��N7@5�J����M䩎#�ߑڧh�{�����CΕ��h�p�sE��6��eܫFEG�F�N�IXqBfH�b������0�$D)�f/�icۓ�*n���<�i�ʄ�e�%�[*Il�N�e�R��d�6�!YȔ�o����N�5F��!Ϻi�`�n�6ԋO��G��}��"�E�K�\a�#>�7�)�:�B";�,�_�*u���k�̎twV��
Mzq��@��D,s=�������i+m\yɅ�m{�>�̟��<s��C��elם�s��>�l��	|��ﳐ5_�SUMPF�:�ټ����P='/X��S�������Y����ɩ�}v�<�!AF����#\	��
N�CAJ٦�/�,"�ĨF��Q��=���N�&%7C`���?��{ơԎËyX���ʓou8)Wґ��⡳\�"^��W�����F�Eٌ`����r�ZP�]����a�WM+�s�&�vǒ�p)BLg�������\���4�qV�JwyR�{<^��/�t�$��L�x���������`q�q�n�_��Gj�q�H����KAP�$>T�P{O��d�o>�l���?e���z�c ����n�����1ut��#����;�u�{������2`�Ϟ?:��ۥ�Tf�`m�NE�8ǲ�Ѓ�O�F :E���z3�f���N�L���Ե��W_����D�},$�#M�K�{�uf��]~��7@4j��Qmc�,����)%�0��q����BsP��B�18���נ��'ʀ����'
&6>@���ǴpL�2S����m9^����2��6*�5�w���U:֋����B''���[�8�4t��&,6>��Zd����8�Hh�ո4sl4�ǯ��BY)"�&Ŀ�nYM :�;��w����^�G�jKt=e��kY����W�Mw�g�I���y�������&���F���4O @z�/�t���߉�x>���)Q�����j�c��-�[�(����Ldv��3*Cnm�@�6�M�:�PIx���Y����	�%���D�K������@)-�j�"t��Il�;��?�S~xe�ՏcP�s �� �p�DӲ�z,]@��~|���xT��'q�NFU�^x��fJu�0�f����~O{��D��`}Y����O���1�se��T8x.���T`Ӫq.܅�� ,����Ы� �!aĮ�� �2_lN���'��6�ǦJ�oc��AL&�b��A��9��� AE��fR�Ѕ�$�#I{��7��"���p����קh�o��R�-q2�q�-�O��[y&�g��mM3J����u���>7ً',!���[ �6�����k�C>�_o��X�|ҞIܔ
Tά�`���)m��ng�����oC<�숦�"l��<m?�M����5����s'߇��׽��+���R�Tx�Kz�4�S�Vx4�ڷ��(�ZD�J��"�#�+UC�(��y��ٺ6Y8�Q�����kH���.l"�#~����5dGC�ڕ.�8�ϑ&���V��S^j�p
V�>s��*Z6�Q�T���r��Q���d����'Y( 4B��,�W��uʗ~n�J��T�A'�&�5��	���˫����Zufѣf���E��UB ӤX�.ؐw\�,1��K�96�BJ%�h�i�£�[��2[��I,HҺ^�a��Wl#�V�����z>x��gN.��R�fH%�8*��G`����Ѻ�����x�7��xp�?)ȁ踮�nm�$��<����36���ǐ��h�h��x��!�@��x�Ǒ9i��햢{�f�]�p�6�`V��ˤ`n󥒩�)̤��*���I]��Q�߆e�UqEU��w}<���j~%a�������}r"��]o�Ǯ&zV'.�ܻ���ߞw�C��M]�%7��.��<o&�FA��x��I��H8�� q��Pܐ���% �%�Ku�T���'7i���D�[W��e���q(�@Y�W���6��ǄI�����1�9�:�^U�W_0v���}`{ً�7m1�w������aF��pD�t0}"dʗclu\F�����!'$߸7������iL��yY����SH�ս�~c\�����W���)����8�%ݳ�N�6�<0�䈔�C�_d��+흪�]�m��G�>܈�������B�7R�ﰅ6>ޫG����k?�
hYp��b�Q��g�>etJUX������{�(v�3�*������r��@���a�i��Aqʨp.|��5��47&���_a�Vՙ��A�����,;U�~~7ޗGi����<>x9B9X�2�E���E�Y⪿�V�"�a42d��h�bIn%#�|s$�$NQAHI����P�7�ͽ�g�@�E��%p��P�j��������_yF*r��n��Zk�Iw�H�T<YR��Cq�z����h�Ä3�4���,­]3��P�2o�r��\3�YFV�S��Nz�
8����L{�r(�l��dHfδ�����Ӱ���@٨�T5lzo��5��rNh󲳖�Qp�fr	˜'��Ed�Gv*�6�2�n��R�̤L7x��K���i�:^~4V��y��Zt�\~V�ڧ��Ya����枿?q�J�����W{m]6hѤ3гZ�����n���c	�5���(�-e��e!��)%�x�x�.�:����>��nǽ��G@/c^Tp��,itw� �9.�C����A�`C���!�x%��_�DeX�̙�`��:/\b���P/a��GY��Q�d�[gl5������ �{��m�i�����B�����B�}����j��R_{�4q�U�ٔ�~o'�����2�ɲ���ݣ��Z�<˥�ON!��"}�i�5ifU�1�@�<W����ª��b0I���s��ւy5)�,"�?�,:�T�v��y9'�3:j��������sS�I)�\�#	�D���vBH��P"P�h�{��5�~,��js��"�+/W^��;e�qq���Ԕ��� �u%�+]<5��[���zN�R� J�LN6�n���jF�r=Ы�DF�k���T�G͝z(w1��
�|a��s�u�=]8���1�<��^�	����T���#�9�x �3��"��K�"|����te7^�nz���~�2��<9��`Y�`_0�9�$��¯����!5��Rn����(ӱ.S�*��>u��g��]�Ǵ��(����dO��bA�c���?���WŬV�q�F����S�W��ps��l�w�~RS;o������bt�g�YW�Ⱦ��|��ڴ�f/��7�c&�F�og���B�.�[� <K��fU��3�|���YG��d�z�+�$/o����q;�AT"���wKR�t{��`U)�e�t!�<��(�lL�\\��"p�����#=�w����wk?�0�0�'�����{3KJ���¹�h3���o�r}`o؉Y���v�P,/����ˎ�V(4���R�ވ�?;��(4������b}Kh���g�ס���F���m��m�IA:����̿����xM�U�3컅c��aGQ�RrF|�����BM�
��ז;�	2�'.Y9�˳�C�#�z�خ�����QZǒv��Z�o�,b�D7�pu��zF�� ��x{�0ϋWe������9�0�X9�w�x�|t�V����K�\ϖ�G�^;�؅#RhLB��P�ɂ��T��ɖ���Xs��n�����3��)}{���-7tу��>�`���b�r������ϱ'�JZ�A�ۂ�,�)M�Կ�E�Tю��G���R�Amſ�Lr���CM��)��}6釐J:����<��`�j�!"ؖɎ����EW�����	�Rm@�
W��K�O�����c��O��iD_0��ܝ����7�IHg����i!�����n�b�dq����]Q��N))o��>r^g/l��[�y=zYm��yٍi�'� <Տ����?�c`ay�I4.����e� VO�݋�f�p�C��;�|o�a�X�x�d~��NK*K��h�[�1gEe(����#��'�D�zԻ�c[�n�%S�__�Ӫs�sH���L�8"ph����uz/�j�C�Q�F��͡���]-tk>������ea���N!��#� �x�- ������N�n=/{i<�)�]F��_���g_K��ְqkx�1�+a|���I�<͔��d���RfA�7�pW�?�$��MWf$1T��t+lOFU�ˬ�BȖ����;g�Ê�v�j+����y�&�S*�%�"~��gQ��Q���[K�"��FR�JX���GISgöw�%����^-��2XJ��?p�y��E�}>��	�=Ǯ�ZZ2*L�o�)�iWQ��Ss�Zq�G����{�	Qj�v��v%�9V5��8Y��4.Bc��Y�� :�[�{���Zst�og&�̫���9��J2�7�V��
j|���޸ɍ��
�+h�S�ŪFZ���~�(�|�a>�� ������)�ςu�s~�gW��j]�bpy�� /�&��xf�.:�HŘ��b�l�;9E�*���w�N_�� hF���D@�P�[��b!dw��\�J��V�
�~^dk�.�+����UB��y��3d�X��c��cpj�{�fU�Ѣ�d�E�ȵ^�	�ƸQJ�Fk��DFAT�7^�N���g�;nܒɃVO�%ri>�$S�lVU0�}ܓ�+~��/���'F���ay��;�AwP|��K s���:����N��	��4��!X<_��p�Ѕ�~��:K���M��k�jw�&B��RT�Uq�N�i�
�Oq8��<hBu�1K���8T��5͢d�W��\k�<�d��Fqt�	v0<f����#��M�*:�d���_l��sBpbǒϪ���FU�塚eE�%j������,�:���F^��E,4�Bj����W��X�ͦ��A��1�����<���E�N�O� �k��-��P�g����R����v�N'���Y���&"a��P�U���E[q�A]�qN��tf@�	)�_b|Q��nm}�>TڑX,G�#N{,�u����T?��-���z�9�R8[��p�2�J��gqҬ�M�MG�2���jz����%�&#p:es(4/��F�{Gw��`���,x��H�:m�h�_�U���V��o�['�+��_bc�����l�3��!r���Aq��|�.i����Ң�I�d���~υ��s�w�� �f���k��!�%.	�;D@Q�'i^tW��(D0���
����Z?/R#8�Z��5|��Q�����PC�״7{��+� I��H�^m������s��9��X�"���?Ax-����Sa4��C�zV�%�e��@M�{'V�Q�����V�b��})H���-Ms��kw�-ȴ��jZ)i�cK����;�̆�8�&���kK�ٛ�8���A���I
�g�m/e�M�'�d^��I>�L�Ѵ~YzfI9�y�1aTׇ�Kbv��l�oŤ
���@�
ɚ�e��(󘧔��7/8
�ppRBRRL4j���~��/tT�X�x� k@�����m���ű����)r�A'�D�P����l*9Ûm�&���q$�����ð[�h��	d�W8�U�5x8m뽷�}x�׿#,��G �X)�IcQ��G����O�U�IϚ���7<;�|Ԑ�Go���J��v{�@=�� �R��pR�Y�W;φc�娌%����e��*|�!�7�~wM�˩
��W�c C�ƭdr�b������f�|X�q�r�� �0�]Q�&��#�
����)���9���=�w2�Sl_W�D0��&$<*�+�̋�x��C�bL��b��b����-�'"�sT���_;+�wމM�]�rRܤН����u0��#��	G8�.�	w�Lr����mN�H��K�d���|�-�%Te�)�r���O���Y]��;�[rx�
�Ҵ��1�پ����-{���E�9@��][W�̸�����RZS�t̮�c�1H�K��m��2�h\VEeK���S��r����tJ����I�$��B�J�d�F���ɞ� ZiP��~{W`a�˖#�EV��d��@5�`��=p�MW[��I��~P�TQ�=�ݙK;=�i[$=�-pqn��U=ۚ"�����O;~y�#�p�;�z	]�`��NPH=���.�l�d��ʲ���v�b�i2�-�I{rԌ�'���g�|6Uq�)�����?��;��:�n����H�G��i�������0���w�t޹�g���Ѡ�k�� z��V���ǖ</��F��s���*��� �l~E>��XC������ɮ�B;9�7�E�?��:h�#�ݚ��hօ��W�����)8~���F��|����Lf����uzZ,t��O����9w�D���f��Z$5榼���>�A��Oa0�U�wFC�8�����Bin0`��=�_T"��+h�ap���K�G�y%IBw���U���s�+_i�єm���4��\����79��:^}Q��I��{O�J�S=n���Q`�I�O`�� {w�Tq����=*n8�/Η��a���ʩ���qk'��}�mR*�`�8Q�!K�ܲɆH{y��ź���6mh���8SD��t��@���<C����@zi�"�)�}��SW�.�%�Y7�Q�j��":O������M�p��Q��
�������~�u^��y8����[DB�	��=H�כz�~5؃�a��*���F��w$�X�_�P�|�X�����J�R+v���'�� Z�/��|>����b�BVU�����G��^O>��>-�v	�r�NF��hO��0��1�-&�6Խ�_�K����ճ���O �Ȏ�We,͖)�TL1��y�������ٟyL�η��(��«����`�c�`k��r���U�}��9Υ��ݶ/R6�`r���&@0J PhٯL ��{ľ�#}D���� {��ɂ�:_�Hp��P�&��CEtJ��{dOd�jn,C�H���;�	���N1��Ϟz���e�2B����5o8�zul�:VI��v(D*��<����������k-2Q�*�5$&*����N�̲-�y֢Vܬl|U"���{d3=c\��6�
D��m��I�m�dH�:� I7y|l	���zI'��?��W�:�L4I��-z 6�)�f8�҄&�6���%�I���S�/��)�D=�}������Da�켉ZoZs���\���N���Q��u��� ��(#��ggQH��ky�U+�$T�&v�O	�̈D���+xG,�����Mez�w�� �qZjk[�k�3{��m~#�PwK˗�T����.�U���O�O��r��|y�v�T��Kԣ�uFD{G�S��5\qd���<c/5��1�Ƕ�H��Ap<s��vثI_.j����N;�?�����#v�E�t?��˲�5;C�ra�� ��.?4�3�U�p�g�$����9����0���p/ 2�������%WHg��'8<;z�͚$-�O�*�c����#Kp�(UV�F�{���5T���^s�ހp1�5��ҿT���1��zևD8��xF���{��Bd�yrAT�Y�ɲ�+i�-P�l�9��F㲬Ӗ{����<�{���m���m��Ք�,�� ��d��r�@�Ε>zʶ��t����&PH5��o,�,FL�
����\�����nM��]Iq0�ո��-��J&x�'\)��(��	4�>��y*:���1I PZ]
����d���=��4�r�Op�W���L�ٯUǫ�oh�ɵ5�i.cL'
c�zq�|�����:�~��u�l�/���
h��[���@�������&,����|�h#��X�Ȕ[�y���0���������U)U: U;��y��3l1]�.�i����S�s�:n��Z�޷UV�=���P*)����!N�V�]�|�*D^T�$v�!���e�߂�{2��z�2JC�����R������v��(&1}�1j.�i�}P ��:৘$�kWs�P���q��6�Ԗ䴚�	n��䭜�[s[�&���E�x$6Ao=���)Hz<����_kZ��p�]��_ޭV�=i�I�g� 'H�M6���^���e���=3�P���Fz����Dr|�tr�L{ �1ȩc`��a��2��H�O�1n��L��&dԝ�������"s�L	�#��)6!ū����+a̯YR܂d�a�93�Ek3R���+o��&޲PjL"�-c�-�.[.9�Xa�N�u�[�u��'�k��yJ��GVp��� ���P`�a�I ����$�mp�~�eP8C�\ҩn�&^)�wi��\�1�f&�b�a���L��T*���#�"�?�w��ڪ���g8/�`������t�oXZ>;�0rXX2x�� c/	�u:%*E3����p��1!�t=^4�6���j�W�<|����.CNBi��3�;�z��ڰ��6�/��Q�zt�Ğ�����������z�oC��H\�'�_�oTSg���P�m�u\���+���̙�K�Ti8)��a?T�8��M�"D�?P6�y�ݴ�,b1� ��Mw�d,�*>�g}4���)���We�k�C�4��L��n�7	~lh�yX\bj��B�Ǆ )���|ES3�c5�2-��E���B6S��7�D�/���p�Jq�S�F�<��bS��'YGL�Rؗ dd������i�a�#SL���g�]�e*�>��KG����SU_�r�$�C�cMvxX�D���3*���?�{�_�~[���_9GX_�x~�>���ԑ�]�d�H8A]���l�_���͎W�����O6�Z��rl�l*��ܠ��V�}��c�5D1���'��&?cZDO�𳚆*�7G}G��-�
}!3G3�'!�T���z����=���ĝm�b��U��N'8tvd����3c��z>;��95����㿃�X>�V�/i3���܂�-]���ZQ��� |h�Qz��-���`�(���G�&�=d�	��X85��@�����SbF��,�������O�N5�OW���M�%\���d��VԭT��T�MQ�<�U�ܼ����EiM}�AD�}&�����!M�32d�鸄��ҭ�%y�;�CD�8gAИ�r�oU�7P�w��R�6@v`@����(���ٴ'����\�|s�aqZ��F��fbO$??�+�#���b��n&�!���jUF�=�����zGK�~��q�T%� yw"�?�T`@�"��͸2��K���@7��Gl��2�� .ƥdJ�p�k|�����_Q�K�Ox��9@7:iAe-zHw0*(p|����鿈X��!&�-�����]���\�*�4����ޣ�Q�5y��B Q$֥]����}O��b
)2�%q6�����ɧH�t�q�m�E4%b�7|�?�~�c�t"%�{�i�˔t�H�R$n�w�XL���p{��ʼ���ey	7u�w3�簳�UkB�q���i�mqF�]�w��a�tG��w��F�֝9��cN7v��$��k���TA��8��O?�v&~hgɠb�-�s��,�1����π1�U�� ��l����n�z�;+4���"�(����0o$R8�Ij>����X���6�}?qBp^�g�/d$��[^n59��S�)���w���Mƴ�P�������nh7�%j�Z_�)@�E���V�ǩ.��	��Z�:��ۊ~g�E{��JUl� &��]�����`T>m�.�N�*�U�9���k_�s����=V�w*/�>��|�aX&,{���J~���Vޅ|�U��E��H�1���v���=Zz\������zU���}�5��&�i][��q����ݔ�D�	影kۤ:�Z�('� ?��]b�-��,�o@`�p�#A
�0��`yq�����!X�&���WZ|<g�k �����A&���J�����'[�Țf����5+^7rk�xD��A�aJ���kj��T^���E���'���g�L��A��`�#��?���~V����1��D��Uſ����~����R�o�3�R��n�ig�-8@�N""�K�o��qH)b��f���{A4�EB��e%g�4֡��(���t���p1�3%/�����m�@{���b˪m{�`N�}K|~ ԉ�T��m)�=.3R��X�Q%�WDN\Q5�̗�Y[ʌ����fC�����$&ù ϋg��Dw~h,��Я|Ȟ9�E�����#�8l�ۀ��8q�V���(C����#��u�HW�⳻EN�g��(v���_��7�1*-������o4�%�_��.ˀZ�r?+l��ҫ�.����x�6��^ʜf,�ߨ>����H4����^�4�����k�z��ȘDI����^�S�i��a����!����Z�w]���U��&����s{�x�}���oSR��Mh��s����ْ���qV�G5�p1t 7*|�Pa�����І8�@�i$���3!΂�I��z�dB+`��4�~_�l�
p�n��}t�=E�:HlԶ)�K{p}���O��ZB3�"��[��KL�ӷ�c�ed�rN�k2m��Ey����h����x��T�g���5�N���t��J�ǁ����^/Zj0V�C��b���ǎv�d�?]��#�NI��9�Ca��#-�����80����OsI0�$����{�NvQj$�\�����"����dV�YIPަ��y�j���O����c:�(ˁ�lKi���܌��Q4�g���cU�z�z�d���l��^�Hs�*�R���
��?��c� �<R��f�0����-�?�=���`L���[�ٲ��L� 3,8��s�o�dqk����,$�&f�̆?��úAxwM�����i���׼�a�*�_u(H,,a]����-M ���xnU`�|۱�M������%���f����(k����[����1�87vh���8G�������~(�(>.�Hk��n`T~,�,X�9q�"\*5� 4�k
�qm�l��
~5�Rk_30��x]k��5=\��WG�	�폽J�^��aF�Ԧ������@�K��"٢��1�nV*<c��b� ��kT�׬D���j"�!�[��N�/�2G�j�o�2��=��Do4`��#���u�Đ	9�n�X��J��/h>� ��և0�g=Y����o/L�����c6C�;�<�d./��Z�������m_�4k�L�Y�8��{�����A���(��t�̺��s���P��r��]$�}�]���t}��w���M'L����OPY,ч{fKf��Z�3VDJ���Ag������c@ٷxjp8W��N�_�#A�L�.j�������)W8��B_sJh|�N�s��v\y��7��K>Rs�F�f�����i(�����d���+��<^g,��U�`����ؖ��R�E*	��Cdm��Z�~�|M�G�B|���)��(�����H�449�IM�tF�5��PB@����He�r�{�m�9�1<��8�Z�A��tp6+�P)���q�M��.�b��+���I�4���e��p~^�p�nnI��^8�}�p��"-U��D룴�"��YJ}s	@���0����E5M�9��؏=V���ڿ#�
 ;��9:��I�*<��w���}��qQ��^v�=�eB�V%����jr���k����'8b�i
HN�t>N�Z��'�4��z�7�v!{�"+c�B1��N��H|T3Yl�������z.w`{�2G�*�p0����i�d��u�אM�,Z��?�N)~/@���	%-��J��R�.�4��_��s [/��3gzi�����Ii9ƽ8A����3jLc_wq�nH����G��x�q�FM������ɿt������j�
�"�A]�9 +^8d۷7e�'�` �KN�
��mJ��01��Mfm��v����F�R�2�02^V��3a�ژ1KI�s�frD�9���Ma���%)3Dh�z3�g�L�Yu����k+
���Y�N�>�WG �b���ϋ���Z���.��$]=R�f�EV����z�]�4�}6�q�&�h6��k��pÄ�׹]9��{���wn�r\�Q�ȦS�6�tt��b{ft�f����̧�u�"�n����잨]�	�8�:��ީ�,�U����?댝�������nG��j,�����H-;�3�Rc����F�rٕ1̻����h�E��W9=�td�����
�s�3Fy�d\tn{��d?��=�j�{��F�6yxj�q/���b�-�K�u�ͮ�+k�j�G�q3��G�i�Cx@\u#��q/�����rϮ4��3>��}���oa������j;}����9�T�W��ΔJ!��ǌTXX9j��H(�Q[�IK[[�虋�u/ӹ����ֶ��!�y�]J�Po��W���9��OIx�1h�h5�9�d�>Q��_=��W�c�5$fEb��I|x����n#*�bz��s*�R�C�!pf�C�4=�š����/�oX�.J/k���؞"����ef�2����(�����͵�����6�����`Ǎ�FY��<�j�}ֵ�6���H��N���D�+H(��К�zcf�x���2 h�yq�����L��O�|���32�G1C�W�Ƞ�_Ux�F�6�����{�`6C�XF0��(�|�� \;H�p�i3�����؂���%w�d���V8�"�r�#'��C��Z�=ìvW�����X� `�D��ޭ��uOȻБhu��Y��i)(`�6��ȵܼ�>	"��f�aY�Hd�>� 쎲�I+s�7��':���V.8�wlv����c�[zY?�S�	�"E�,����c����*a�؞!LL��8_3^�t3����]������o��%��uOS����{'�:��I1�`�p�OkH*~�:bՄ��{.�Iu�pd��V�[iԥ������R;�4�\C$p9h��-����O��3���ZSB���@��xN�1� �� ����-�(�O�ҡ�=j�j�b��P��gQ�*l��F~�ʇ��&��H�ǒ��g�ԡ{��G�l%�{4�ߥ&E H�k;�w�\�^�b%J�c�r�{]����ZT���&��,>�����a�����|g��q�������<hc�d֠n`����	�=�"\�h ��H} �3�U��:h�se��&:��h������ȭѴ�p�r���~"�T6��C�b�H���HY��I�S��J�x����Gt�?^nƌ!Ԑ,֡VZpV;���~\<�3��y�$%�GD�隣��y�	��5��!��q+�;��ٙ2L`X^�B�w��HI��W���ە'��}§�K��X�\��cT4��yʕ7�g��
Ӎ�.��%-��W��l�a� q�6P	vrKl����_�mZ*����q����~{��0�@��I��ȾK��� ��́)3r�Ѥ������;��|��D h�����@�]��K�6Bp`m�qzq���� yr�.��~�[�<���t[� �6������_}�}���u
6KS�Nl
��Q+m8�z̋�Qܪ���!��M	�K�r��*��C\�&Cr&�ҐA*��W;W����_�N��~����.᷎]�g��GL�P��*Ec,J���'�B���7"�xn����xf��~�=���o�a�(�Uճ�g|��`�P��s��Ꙁ�zi�re�0D�����$9jN�bk-
�>� [۟u]p]-0�z�/�[�{��b��>����@�W ��ǅ�� S��I���}$rLR�o3�lȎ/��0��σ��kBD��	oщ�{�!L�'>���.�a��
�7��i���:��N���w��0#g�k\���ޱT0V�QGڗ��R%�kNp�uO{�'vl���ɐR����;�w_��DZ�y�t�ЖtDqN�0�����3��ڌtަ������X�ϕ.$�&J�����a�����q.��@�RG�-��� �e�=L���\G�qrQ�� �ꍂ���z��,A0W)��9SV;0�? �mI|���W����}�1D�q�hW�WE�=��eÂwY��(N!R���S���My�j�?B8,�˾������/f�(�aov���ؑC�W78-�9Q�ި��*}2�L|���ct�SЀ���w��>F=���D��q�c�����4�v�<9�.�S�����Ð���%�h�\ƞWF��g6 �p�a�/�5I��L���𤌃��ߺi �uW��v�����1����w1��7l�a"}��dx<��uzj�@��I,'���2�$�!jF�.�Ⱦq�(��V�2?x��ñXχ�_���k]�6h�MeY<�=�P�\RІ�j���(�z���W�difyl5O�B4��M�r��D)���T��Bk�x��>M��C�^��i�U\�8�`bm�ΈX�o0�X�z�Zt�w���,9�-0�8��Sし3;GJ8U�=@>��
�Y�9�Ɋ?Qd����>�[��3�-m�0d.�[�@�UU6���k0�S���ò��!����(����$.���(:���Y����{V��&=yF�TK����e���
N�4�π~n#���!h��x\f������=������g�ʹ�����2ܮp$��W�u���; Ŋ���a��k|aڹ���m;��(�ĠxiT垓���_�r��V��2��<�UCp�<J6js�i�ظ��3N	L4�z2�6np���1��[T圳s�M�������Ɯ�d<�
w�?�d�0�w��ʎ�C.��}R��h�����mSkE_
�ދ;�Zp����kP�#�l_����[�%kf�I,�r���kЯb�i�AH��*G���^l����#�DCԕ-k3{�F#"�k9YV�B˦�o��K#���'Znn�Q�AE"ٞQ��5�u'�`6���"�	���̴�|[>�!ȇ��h��s2SC�g��/�+x sxʨ��F�GWlR^c$z��Q>���u1bQ���;�O#���w��S��v\m~�펷�V���D�Y]� b�������pN�����xp�˩�D�فZ��׶���I�D�P�d1XX���}G���R1= ��_��pj��������*@b���W�o�U]{���\��`��Q<[r�-��Φ�K�i�=�O3f��R@�>y����Y�:p#����ڬ簅��8��㬣�n�8�-�2�C{��QZ7�ʦ��FJBjL1'V-i�u�~�K��	�<�>����ğ��5�=��k_6��<f�uB�9�.�;O��n���؜%-���cÂb|t��O\6,8*wj��umGV#�!vę�!�\��S-Fs�9̶:���#��������5O�(�2���d�z�,-���y���۹������7nFd|�`��y���x�.�y�ί�0�!��S�v�X�G�rOF��	o���v�jPk����J�s��\��Ç��������K,:4@�9�~�F�0WC�Ωo(��D����G9���5g��ؖ)�2&x�Y��ބӇ�Bi�n3aP1Q�w�%�a/_b%��-S�ܠ��i�ٸih�: ����`��a��"�qp  ��ˆJn�rL���=�G�/��~���y��$`>�� � ��)��b�MG�!P�cbU$2Ȅ1�:J��決�w�  $�����	�۴&����#�'�^n�?�5Nlc���󁫭�>�*{n�k���|�q��`.��.����R��s��f�2�&�\���WPl[cq�i}xj5��l��V��e���-�	bTU��t��83}�q ���KnK<@q����拺a��AuW��-~ A�<�Fе�x�%�V���I|�8��qO|�������ja�׿�k�_�T��h�ϗ�d�E&�lX��$��V[W)�� �x�-,��z��ڠ��cTV+�Q����䚺�T�,� 5�� j��ˆ4��U�N��	�_+7�N̳�7�ZN�wɱ���3���ֆH����V\�bY�!��:��ȧibd������1����`��v�<�̛�M�LQ7�g�Y���k�����ט'�U�߹4����x�{��n��sA}�b�#�t~,������	;GNh]�>�d�ɡ��[�܅u	��Z�ʯO�h����Bb(�n����#����$<�J�n�PI�@��ݲa�`ڧ�6,%{
©q��œz���P�/���$�n��.I�)+�A��M���[�j��	�0W���� ���pz���tK���TKyc*�Q�KE����υ�|��0`e�]y���ZS!&�hz���&-����-��;�0�e-B3H/��;rr%��������\�$؅�+��$�$_�+e�bC�����	<OԆ$V.�ub
�Ov{�/FT��w2Sk|<���%A���F/p�|B�4��*����Y(�*��6t՘n��}ݟ=���8�*��
����Y�3�k��U��s�p����d �4�(cI��E�ZV����r�`'m>�t!\��E���2݆�+ͅ���G�U#s��;�`d�QT!�T���{�m�^.4P�*��Ak�ܪ��*��c�6�9�
���G��r>V]�1u��pv���f;��e�(.f8��i���ޞ�Ox�����SوF�D[R��Loj�qC��-��P� �9Yb���r��0�!�&��e�{��!����!JX��؟��s��}����T֜�R��ls݆�k��0��.��ڼQ $�P�ԓ�g����q�π�{vh�?��Nv��w�~1��`�`�*HQ(�^�e�j��~5��=a��a�Y�#9ǎ+�9�y�CB�r��{>�ƻ(��24�㐑����	��Vi���� 
�$�ۖ�5��T�@?3L��b����'�R"[g��V	�)D(X��s�Zb!��`���w��Bɵ~�<S`V|���4�uq����Eʅ����IQu�x��Hy�,n*��Y�أ��:�V����V��F�"������07����`���ա�����@���̒5͑+�p��hS���BDQ�-�:P�C��v��?P��,�a�Az棥n�����B�0�fܖ�/S�M2�o
[xzg�[�"����]�ꦫ෥\^��D_�0��2����wvdo8#T_6�M�jYxB�yT5���$��:N��a�@*��2��_-�ŗ�P��:�����&�,�� �Ҙ툉�\����ۅ������r�@��%�g�����=f�>�t�6���ANZ~����B=���6o��l�f���A��>:��@�9�4��5][k�ҝ��tD8���d�;~�@r�����Q �@N�n�4�u�>2�'$����7cm>J�S;�W���ǡ�s�H����~]������9��l޹0�Q�2i_�_Y/bl�ݸ(j�݌���!�Qc}��%����<~n����Aw�Q�X��m!�c܏���$TAs�@� �A��"W�`�oc)�c�Tȧ�luj�4��S#^���y`(��m�f�`W_)P�9ŵ��'���n ���K;N�>&ZÆ�S�N�܎g�y ;�F�\�W]��	��6Sy'˪Vg3�u�x��A�y8-P�\a�ny���q�w"4i}|��_�}����2�g���w�L1=h߹nud�{'`����1���H���p�a����(c�	ρ�m^6�,#x�4�_�^��:b�7�t��t�S�XOA�ֿ�����c�|k�bY��Z�pA���C. .}�ے��BSŔ&�YI�Ꙭ �)?%��9+'K���d�&�@��D��}�I)�#m�3U�%�bwn&��+���{�_q���k`����'3]���ۍ�`��
��=�V��1��\ڲAqZ�'}�����b#���{6g�����"olJ��Q�<� !0��(%1o�,J~�`���0���Z\Q��6edX�Eh�4�$e `���M�����w)=<?J\��ET��aM>|�~�?�=��в�����&$E��rU0RUə�)�����
�9�QѠ�I�N�.�pN�������p����2��Ig!\�6���a����r��Z��tr��eW�p�~���%�i�ws��U�/�I;�+����$�g�IBU�m�!��%����5�o�b�qyn��!/u����.�#QX>��ׂ{(��A�`��,�$O���� ��E�y�RS\�F6O�Luk�D3wVh�*�r������b��qքz�9S;If��zF/��'�ݺ�p�F9�NA��.Q�N�I�vD}��oe8��C���J(��v�ҴY��p�X���I��
�Ue>�� YU�p�U~�g�j�N7��m���޿��6��Dh����­��f������@�C{�w�p���^}���3���6'�W��������[�%�l�e�/k�x[��>��M0#(�e���p��t$�6���#���Jo|�T��m[�u�}��Ui�j&��Q�\_�M`�*���6�
ï�=!�9�;�(�5�g�ޏ��REpˆu�q�O������� wq��z�#�X dt{�-���x ՙ���c���@�*[,��k�b}:k����+."�7(�2ʽ[J�v9X`���:%��Y���Ј#¤�.�M�ؙ��x�=盱�3H�N
���$G/'ǹ��|R��	wt&4-%��4a�DcFhx�8���}^^eF$D����v>�k���$l/�Q_>� �ՎVJ��o�"�3�
���2Y{���=\| >E��iP>� ����[�H����U��
�}�q" I���*��&u)h�u��ulm�(��Vo+}臬x��h�KsSRL~��+�_�*"�Yqk����k�1����n�͊8�WJl��
't%�����2��d��e�5���`�G��[����,s�,@e#ܱ�Qt&��?ƙ/΢@�R��6-�Ip�L"'UIs�LO>�rGu��3���ot�\~��_�de�k�K0�G�m;�����ړ5ٖo�E!�P":�߯��p�9A�@���sV�4u�7J����)����n-�o�������gJ'Z��G�aMٌ���[��Q�u_$��k�b�ar�����q���w�Ek���V$O�.�&n��3���}%.���q5�?z�C�_�?��RV�\���aAH��,�������2뮏NU�
� k_+S��3Ųb��OX��u½�E�$9�D>�z'��1�#��� }*sQ�����(|���6����^[��A��}�}'�q�o��kl�{�2���Ej?\��n��`����	��񲥎x6��(������� ���L�A�eu$�������)�o�>������S�Ȕ.�]�-�B9��U�B�y$��nU=��56q:T�jr0ͿÔ��QmP%�|��r��9���U�!h㪀D$�G�W��9p�E�2D}�k��M�q\`)�5��>e���Qk��ʾ�Y���l���"�'�Z=�fI�)���xe� ��#e��d ��>� l~sҬmQ^��p2Y+�MӅ[��k��!��S�4�*�$���V���6ggl���<�&�,o��a���2���%����{�08
��
b�^���z���@���&�>p�Ώ�ʊ�;��	��ݙ�`��R:%ҷ��+o�D kNXI�'�V�դ�&�իkh�v����K���WG"��`����'[��Y��
��b�>���Nh��ϳ)Z����b��v弶�B&٠����SVj�9�l�����+gD�*��2dcD֮Lk,-���E`�>�8�5��F�v[1P�s��@)G�N�i����O��5�O�De*�����D]F��U3:S�=*��l�Z����'�������x;�=O��L��LEuZw�<�1�f����ӊJs��:���6�d��Fp@�����<U2z�K�zh�7ҥ+�����l�rK2�A���'�r�ķ�e��M9�)�+�H�[�O��8ɣ����^�I`Vͣ���o$]�8���BI��M�JH�wh�o9��ë]%�G��MJ{����q�]�G�"6�yf���7G���_�w�F��Y��y�y��3�\�X��٣m��fx��>��$~Q��`��}�<è��H�_���}�+�c[�Ai\� GDި%Qa.��{� �0����F��f!�]廚���B�ά ��mt��'42�gJ3>�D�Q{Z�JF�zD�J�V�(��@Y�}1�O�����R<	��*�e�C/������X��\��m
��kXs�.˵�w� lx$�W���۳ӫ!u����o�lq:�(���M�r�Ϝs�9�9�pI6��.ʼ��r:s�Bt�&3�.b�c ��m���t �p�����*�.�fCgn-o�����+���7NJ����P�*�>����=��r�ڼ�Rm�;��at��Ō8Q����Q�P&��E��CR"~�ϻ��S�|8����=�|�&�v��[��!�}?��F�,j����?#C�ׂ]�Y �N ii�o�B��9T�\��������x�f'+���?U�2�R�ո�\h�����O�m!�i��3d� �0뗑UO��A3L�k��7k3��n%gQ�����w�=�����a�͖@J���̊�*$LՑ�I��r��,	b�X�y����˛1Z����,PO�����'\���0g�bԯ<��ŏ9�y� ����\66�h�����;��l��7�u�$��ɸ�#I��32R�0u2��,*<�b^�����<����N�a~�`�xM�؜w�X;���	ԇ�ܿ�漬��;���J�P���-�'�c�,�·n�"<�m,�U"���b�� ��\+&
�܁�堔�ks}h+�`����67��;/���!=�'���|E�(���%��+W%,���J���IXO��}��o��YT�o�ܤ�q�f��/�K�E��'n�qrS�{��{�	�8���=�{�����2���q��X�P�vg>�UW�ֿ�H�d�N��Cʝ� �D>�.��D�p� Y�B;��H��ʀ9��Y6i�Dn��,$�^�Y{5��^�!G�:9���KDîO�X���� �����o�1�:�C�]�Z4l~��!]�Ll� �������L����Q�##�,ٻv�X��wP��ZZ8ē��L1���\*R�E~��h�":��{��w�&��/�P}pko�V~7Dc�'\���d�ꟓ�(6}"����au�|Y�	x^\�.?aDӌ��Q%\o�M�¾ɟO��h��}X��X �3��.q�S�S��G���_��;]��|\&�9ѵ�A�e�I5\a
�/�ؑT}k�x@cb�}l��bz��0b�:-u�w��)��qT��Lۡh��0�GΏ�Qt��j
�.��ĮWj���"�SKަ �t���������u��-���w�0~�H;@��r7j��LN'2�f?x�X3�59��s0��5��� x��Zo�\��,�;K�&<NmD���"jCm��<tw��q��-f"i�&��/��h�nI��(�P��v�7�
�(�o�\�5�Չv#!��$H|Ҥ�[Z�T_��-����w?��r�g(M��A!�
g���
�R�#؈�0�-b�� L�r��T��<=���gf{�S�=��a�^�I���������` ��E�(Z�/��;��@E!T�'n
�-���RD��&�ҿ�vW����!��A|��0��ӿ�	�	�C�֚U��A�g��D-l�w�Bt�d-��I1�<���m �䂱TRh���9���ݨ�ɾk7��79�V�CL��\�S����ڨ7����E�0A3��5̦:~N�b��/]�*�;���9�S˓�_�|+q-��g����Cvʖ\`qb�%͈�q�x ?,�@�C:��T�`+G���c�U�!��p'�i�"�9v(П�E��q%�2��N���6Zk;?�W ���4��e�faA`u�R�m��15;��ڱ�T�+�����DӨ������������ʵ_��f{�!�<�x�-�l�c}#�M
T)�+����~%�xy����4C�G�P��M�Q/&^Ϣ��ͧ_Z�`����>���[�ۜ����R��a��KD�E��| ���ݔu�qi�O�$�\0O8He�pG��Z���x��8g�&n�b���4C���r"�S�(߽�~DN5�>�.B���6`�௬y���׮
0�A %��a]t�hy�fY���7�����u�h ��J�+�RTzR�
��"0g�[���n5��R�xFS��	R������3,�⴮�* T��OQK�|����FD��^��,@9���B������S÷Df�C�t3��5O��_�8k�c5K;��~���@�v�1T���
c����Y�N^#��&	����ȳ.��3��CA����K���j��9BUM[B�:kW�b�r��?L����c7KK�V`�f�^��}	��b�1�>R�\-����GאIz��ME�.S�5���ܷo`u&z:�� N.����0йP�mѮ�Gd�0(����56�� Dϔ�2��s�Fa)PO�W�Vx�`iސ��|
@���Q��Kb'm�c�p�'{���c��,�?�C��S�_�pn�XS?�KOƸK�$Uxp�8[��H�r���T�_��DvJ�qeIJ	@s�u�^���X���To���o��n�A�4�L�ePս}�|k�W�[��1��ĥ5�]�W��զ����JW�P��Ȼ�U����܈Kt)��
�f�Q��;Cq4#ϻ�T��!�>�K�@n��RiM3YL.Q�x��#�#�ZOɷ��,���8v�@
��S��P�!е��Z��$���]��s�`B����䝩Ҍ�P��z������W�v�J�D4����Q3��1kiw�W�|��}=KƌJ����h��<�&��C�V�n�m��T8�	��������(y�sy0�;���c�h�]���Ǡ�%2�F<K�W�8��b��D,M�j�u'�#�K��g)�5y���f��{�8�$��� &��:�ɵu*�5[�~/��bX� jKO�k�U\�E�̱�8�n�n]lQ=�G�
�껠��Yā-7�\Z�y��L��~�Q��p/�6��3��ѷҌ*(nkM��e��		����;kN���.t�'�]��C~k}��&*~���8�"�zU�a��nO�h���B��٘���JNb���1vW��&�7���]�����U�%��'v�#��*˰) Y�G��f��K���Gώ���9L@$�v����u5�!�.�j���
��0�'ב���y G�Ǌ����Wr558�j<��S�n�=�a��#�#2�X��>9�������P�˶�.�r� �&�G�g}sKpE��vp�϶��6�F*%�F�s�	�q*D[���r@{\�О3�d]z���Ӵv�/>>��Yy���wٽ6��qܯ��:6k�H�V01���^��H��gT�m�&��9� �!�~��n%���`�_��)B\���2��X�Q�B�?�@���JM7dnE�*�+M����p1(m�8)|��9�M�:�����ɯMZ��58�$����j�tmo��;�A�f&1@I���F]Vh@�/(!7E\D\�����6ER
5n�J$ap���Z̻w�6����B��q�~�)>�w9Q��cxT�[�������@���J�g~�*$g����V�:W������s��_�R���K��O]�s�X���u)kn��)O�k��I
��6���5�\��n�e2~T���Q�c�k��t�p�'�H�=�����ȗ��ǋJ�X���-��s"dc��v�F	1S4�F��H���Lt��ÊM:*�3GA��_;/���Df�$ӝ�ė��l���^ch�H��ȅ�g��g%iNx����G�_)D��y��������j*\������÷3s8��B��FB�rqĶ�I�lY�¸#�R��Hi��qe���� 8�2���K
�AB��ql��+��ף�Q�?����KT�|~�{�&�!���T4	4}��9�gs����w�1�=iB����'�:�� ^A8�*,Yזb���D���r|��M�,[N9Z� +������(1�D�S�Za�h��	��@�R'�:�H����]�<;9���y=���
ZB�h�&���'�+~#@ǝ�T'�"!fC��{� 4��P=��f��������\
p8+Ӝ���*�.��@v�'��-�0HCty�Jf�|z���h������ȝ^;�U����������g�Cv(��d�C�}�f?�-�hx���7����m�Qz
'Q����9�e��~B��+f�_0�35��]�X&>��˕?��㸜�f�OK�4`A��[y!Wm��&�0�mdf��ݞ�� �u&|?��YM&c���	�SX������6H�O|�5) ��y��Ԇ�������O��,�>���A#�8ve��\43}�����8���P�������:��J*��Ԯ:�����uc�<��g-h$/3�e�w�9��Jvk�,LE����]Db=뻗�X�8����.�1*���+#�u9��i�t�6�pOp̂� J5(���c���ǝ'�����'<cO���O��PE�uH���,���m�Z�M����l��nT'`:.���w��R٨R��4��w�;C�`��^!��??�|��嫁d[/C�I"Q���:�q��X~�d��x�Mĭ�Qbs�P�	3C.���Bi\߄̟%O�=oci�VH��8N��})kv|4�z���o�,|�5�w�Jom"�;���0�2.�t��L[�)
������%V6����02$��뮤Q�hE�P|��y������2���:����������g?��X�0p�I�-A�`� ��5��ei��[S����oı�៖��Hc";l�&]�y�Z>����g�1�^���R��(A?hU��.�
S�=���de#|B3��������Q�1�>�0uLH��Y��1�lk�Y)@g�ȵ��~�y��23m���TYr�ױrz�
 
A5<�K2L@���~�2z�����o1Z���sq������H�D{:܃��iUY��So�k����za|K�gx�'�V�������G־��R�?h��-������}zp�%;;��̯,�]�2�i��%�R}��=zqޞ� �J8�!�X��k5��\��;$�O�Oe��2e����3��m��ob!}w4l�<�����مJ	h�2���-u=ɷ�Y+��4�`1�$#,��3��si���_�'�D`E y�#�p�L���-��x(��̐��8��ۗ�-A5Dc���xc`��x>��\��5�� *^lH��絤��A.x*�<e�{��膩'���5�Hޘb���7:�NŻ�I�S���-�p������|�[�n�W�중�L���,�[���e�:\�����g(J@=k>b����=�XPS�`�3�f�	�1�q&�]�/zt����0�~�Ӏ��ΕQ�V�v�D5�v�o1�%�r̴6$*�
I.��*�f�3T$�y��aH`'ľU��O(��;1��ֹQb]_�s�X�t�q�td��K���M�-d�z��0_hT���i��P�ව՜謓ԅ1�{�:u�cQZDβ5>atR<�����"Z����L���i΋kM�|DyXy�"�-E�4�Iz�xK�Ȼ�r�_��2�P:�ba�ߤ,[��$ra˥ّwA:���3��WS:�5	g}�q�����*X��Ш���x�؉����o~/�G٫��m�/hq�6Q�|L�8;p�����x��?&M��K>¨���}K����|�0�rj��6����⒘hU�1�RRP��t�Oew��:`�f�+��J&*�+_t�!]'!�\�u�sɠrK��$����9��s�ѡ*Xo����i�P���{��RN���QͿ�o���s�+��*���x��d��'�h� :Wd�,�����g����4b9�<a��v��m��/������n�ɶ����Н��Ff����o@9��t� q��P0�˞�'B,���y�"8����ݘѐ���F@F�S�'��&:7�sO�	-ރ/I��`��	���黂�N 2���(Z"DV���1���i�r���~��9EZ#��B������hh��%�5Z���K�ջg��xC�^����#��2��A�Ԥ�Ȝ��&���<�0������U#�f�4ğ�] k�ο�����I�5��mͲ\�n���9��(��P�ӫ�Y~yL����l� ��ځ���wM���l�MM{�ԶXrY(�
�#OEN��^�?�4u�q,�15gñt�@�v�Q���+���<>����F����Q�%��[*���]�Q�j���m���a ��+"
Z$�Fj��Ĉ*����(���%z ��i�?��p0Rx��@G�{|�#�Tn�G�1��e^ф�?LZ�`O�f�tGgh�q/vNW�E��ΒRIt�k���'�`;�2���:]�>Y�Z{�V�Ŀm(��6��Wc����;Ny�P�#5[skpN�-({��+�HYUv!�gwmX�m��g|��m�Y}�b�٥}d~��o(g�~�D��=���r��n��ª�"�}e��Ĉ��k��j����?�A65x�d�ƙ.k�D�`�0Kh�ˡ��<)k�x���ݙ&����V����#�I�# �}"�&d��T�_u�d��N�3�����83:4���8��=�!�Hr}�A쏂�^q�5$؄x8�7��:k�H���(�m�t�!�N��8X2�Af��7�n���A1��X>�����W@�rYm8�@RCը��ټ����%�i+W淀<��o	��#��i���`���]��kO�p�-��{nxƄC�C���\�(�	
4�i _T�b�%bĎ�0��R�Q[����O��I��k#|�7=�MRx�C�̳Z�SP���&n�j��	Ѻ���Lf~>���3�4z���zӹ)qۀ2�˿I�ǹ��=���h`""��hbli���0ԙ��#��۪\��c3�^���D��L�B;n�(h���E'lc�Û]rh�!y~�a��4��U8��W�C��L���b�4��|kt�'=\6%D���4f}r|D#h��B���6�"�����-P�� �_H& 9%�S�{�2���2|����)hڃ��GbG��滻��I��&t�3��.Qo�*�[�U �K�&
�9���Ѫ��2m#GD�A5b��B�*�&�Q�e
�q"�OǺ4����P%������n���l�@r�<�L���2�;-Z����9�*oo]��Q�I��3�m̮��
RsWok���q��	|��}0��ι�������1�v��v�R����3���`����&'� &Yy��U.Ȏ6x&�D7�Xۄ��\��̎B��A�;?�+26|�kb=>�y%W#3�_F�U�c�ien�Z�)�fC�<?L����Wϖ d;K���I�ʌ���K��	O��JJ���"8;|��a8�0����((��}8��̋��`)�v�/]x��#�?	���d��]��a$��� �C��0 �E�
C�6��� �8X[�K@ʬ��,�[ռ���mº6�R�^"�Pb�S���K�q��ő�J^�m �����߻l�Xy#Y~�5Js�����^����"��KP��Hf�iaj�V�7�C[�&�h)���^��\�Kg �����ù��-m&!���D
<O�
�9���!�1����0�8E�/������&1�O i#�p����Y�~wD�z�Eo�8h�Ze}�*9�DK�z������<�tR�8xaH�,- ���E��\���M��Y�����7���71�!�	-�K�W�4i���GFA�R���wM�a&��2���$`~��~�#�rr/��g�A5� :��mQ��H-���$<�<��*�	 �������$�m�Y�o���}���2͠5�;�d��t��䎿��ALe�ݺJ�:&�C�4j:*^�����yG�����l�Zn��C� �ى"��Mנ&�Y���2�\/�gi1 	����M@�/��Q�@-����9�sG�u���9Fט���J�:Mc���ͥRٖ�k��jo�;ⷾ!�����,26@vx㥕t]�ob�>��}06.˓<u{y���vjo.�BH�\ai�;��5kbI����=����Uc�$���O]^�u�`~6Dn�%��;3A�
WӓR�^I�����:�Vz������3\!�jk�|�V	��X7S6�g��"�7��ܻ��Gsj�ۙ[����En9WD��`�ZX���}�~�������:��ߵ�qW�O/ �@��1�u̍ΎV�'0󱜰z�1��ʻ� 6�;H���z���MQ3��i�QH�O� �qu=3�ה���w"�x�.$�1E�K6����`��Nn���0�D��v�6$��g��v�1�h�K<�'��+%G?�O ���ߟ��J�D<*�%��{�:��C�~b=���[���5�����ö�r[& ��W����&R�oR�����(|Щlm�9��;�~�H~�'Έ�L%H)�D�d���HD��ɥ����&&6;�킃X�t;Qn�*���F�i�j�&=�.wY���[��� )���f���:)����vY�or��&�F�O����Au�J�=sb���	8I�R�@�r������[|�4_�O	x*�U�(�~|����rFiMfer+zO�g����,V�4{�u#�n�*5O+oN�/����<͖3���\RJ��x4�OI�M�
Lv�(��o��i�|Y�g%)�b�d�o��r��MT�_�?/N
D��
��>��X��=ׯ݄Y���3�
#��x�%?�������
�_4��/����e�)������3�mc�}�{���"��>B �;@4[\�G�I��"� >�Z�qG�q����I�#��8(��k~�`#GNV��W6[�ƀ���$F�'��uF�:�	�ꦩ����|�aR��JGQ�<�x��F9�U��ܸ���x>p})UΡ_e��t��_�R�:��Yu�䪮�i�|��Y�]�Pv��l��c�~�H���ęD��T}��Ø3!�N�ۖ���	�u�^V|j�g��3�|���0��z�v潊��yɆ�N�n��`��I���s35�5�Nqi�H|�?�X�`pN��«�}m|얻xD�H���}�.Wj+�y����/�(���Z�`D��+c2� �4 ���eRx�9͜�c����0I�������i�|�=��̶��4�+9�ō�:��ilX:)?0�F�#^\2�-�L��vKs��8P0���71��$�kz����kJu�P
��
�͔9ܐ�J�qք��������xe<٨<tŖ�����ʈMȌ�`Q�>��,v��,%ġ;�A������.�N�X�dk�%�i���i�,��5*�m ��^,��_�Fgܩ�/�4�ȡ���_���M�H
֤G��օAe7��]�{�>�ZĹ�&l��G�I�M���+��I~Ç�)��$�c���W�p���u�q�nlNP�h����:eq��0�����O��C��Ʋ���z��H�8S��幣��!3�L��s]�X�D��LV�������Q���xX�V�2�{��$_U�m6�1�O. +���y"��/;��������d����˫c�D�<7<�77l���˧(8$��D�M��Y��'um��*��$�� LC.>����������ئII5���)@L�J}gf�'�s�i��L�x�����}D_r�Vh �X�U#TE6�W�U�5�(5ݳL�_:�?���;1�;*V`!���f]9���|�V�|N�~"Y2���G���E�"Ҭ�QKh�X�j��nx�RVhG$�䥷ϩ�aD�7Q��u5��N�c��W@ y�H^]�}�����@k2�'��R;�t�������w�#j�+y�q�M�/�xIA8�0��h�L��u�׃%O�ѧh-���oS衕`�����l.�T�5Oj$pHY���y_�r��+kz��Z���m:��|[u�K����hV��t���bx��Z <���+�9uϪXXx�+��/J̹v�3�7&��xcK7F%�	��C��Ap��r5U�$��)�+��W���f6;��Z|��{8W�36�s�ݎb�iE3��
KѤ�������{�n*����ڙڔOY�=`�����T���#� ����N��[V�Q�u�k�{o&�þw�V����V�~��7A�^?�<�5��?��>��
���`!���Z�;������}~�8��j=��(��(��˧nH�U����6z*��S���p����x�	;�6����?�K�l�"_�:�&��q�Qi0�zA?��'�Ϸ��	�5�h������Yb�D.��!K)�:.�����	�{�����?��f=$�δ�LME�/�vRޛ<�7� :/�'TlzY�l�?��ʤ.k��~X�	��(��G��ƛ��#NS���)|��H-��p-l�6�5)���)/�k9�W��pY� E�o�����c�W�g'ο?�Z�H	W���v��޵|���2���kOQ�"�׃����ٶ���<-E��n�&�$�D~纶�C��nC�Я�T�j�oр�k",^՚'����c�~�GQ�b�h!)��ֲ��T[�a�yA%�ʖ�c�s4,�_Au�J��'���B\ٗ�OKs!<~YP�m7�p�Ƴ�޴aCS�}��*:�?d�i�"�=��0~n�FD�r��TÀw1b�v��2�<4��D�rڑI���qb�,MQ�u�uZD[^ ����j:yz8(=���0����X�qn��=��M�w ���DpY�C·(�"�Y���C.�A��4˪�3d�c9��cY&FMS�٪rc�34DɆ�l�1��m����Y*�~�h�H��q����YL<�so��{]:jb���ea�k���F�Z�Xv�Jg���K&�T���#�tme�j�h��%B�	U�Ո��	�|U�J����q��k T_���6����hrtCP�J����Q�"�p�$�n��b�f̆���&��M<��>�yg+�����SU4�:�kO�V-\	����PO��J\�0�QTQ��8�"o��80�����/e�xȢ7��-�o���W�Z��}_�hW�LX�dZ��Br{��h1y5GEDt�\��f[ۛY�ф�eЯ���"��$g$?�U���T�pں�1�@�Z�P�8ۗ�-�����+,���"O���
Я����/V��i]bYDmou�m��_�/3�N,�0l��@���6���\�U��xL���[ |���̊��.ң6���E7�e�jr�EB�$i轋laen�LKwV���s尜}ҹ"��h�	iߠ���*�|i�{o���Di��}��B�u,A�X��T��b;�H���z��u�II&+8|������ "o6Vixd8:η}!m��)9�m#��	;�7��M��Y�&�6
��;��ұs��*@�}}V?���f����l�u&[=�!$`�^�����6�v%����_	ou�L�\j�=�^�S���.��.�`!H)f�9�Tw`��@�!j[��7�[��	��� �٪ݠ�X7��2������*���)m�hF�75�ꬰ49����EG;^��2h��\�J~��;*T��,�T����U��ܷ�k�1S1���������
����p��2MYy=�c����t�L�t�D���o�$�E't��� �m̚�d�>�!x�6D$�?Lɭҷ�M���VX�$Ң%��Xڡ�������֛�k��u�T�y�v-�� }1��
/KVx:ɰm�>�9�M��T�ս��>�
��P/y�|�9ܢ�M�i�3����IR�R{T+3Z�@%7��a%�/�F�iҽ�}I�.O��e5
f�WHgeI)d%U���}\��>�͠y��Vel�×b;RJ��_ ���3i�^���˙��aӃ����+��pB��,6�vE?������{��O�_FOӇ���tj~�P��{]�M����l���c}R\ߐd���&$�>� Sw�40�)����U
L4BK�jB[jG�%����@Q��%$�		�)���i�O�aB�v^]fB��,Oct}������i�Z�$/b���l�͡|'R+�+�To�t��]ȡ��	����!{1�8���?�˸K� ���U�B� m�4�=eI(Z(�_����-eB��B�"$��O�۔�.%�]	q2��	]��`3k��ƿ��I�[���@�|�J���
v����PW�ͻ����X[�^�l^M��#O�M���;>!5�+o��"f�+qp<H��Q�C	�T���:�N-g�#�l�t��|��M�t>.��e=�ѳ^n���1�99K+���̲�N�h�$>��:�B��T]M�ԅ��¡����i��TF��!`Q�^&�7��^'܁�Z`�Ջk��c��3>v-O���N"La\'�	�g"9Z�p��?��J��Tr��&j�S#_?ϴ�q ��N7�[��?���NƔ�=T����\��W��֛��t��i���w/�s]���ɧ#7��MD2{�<�&@�S�PL�:���e�~Z /�T�m�,��£0i��I\7VS�� ��U�u}�rzY���M�*��Q�vdlͩ'.�� ��*4FޢY�����5ͩdw�!5�����'n�P��v�	�������񧰌~�ӻ����1utFD��;�`��E��^�5P����z$��I -CBԍdDN�Qq��Ҏ���ê⠂8k��X�m��K�^Ʈ�R/|	Si}ғ	��?'H����|[�U)Օw�u³%����;3=�1$m�3� 4��Wш`���n,���ER�U-�v~NQ���;��X����;V�J�Il]5�r����&�e�Vt�����*�ʮ���	;�8��{��Ҧͱ�'���؅ݱ�#z��)op���;N�؆d�z��bVvSƋ���j���"�-b��ב���������奖Q�e�-�K�U�������O1��
(���s*�������������(�9`��:����,ԁz|>��9�(��O��rj0�d�:Y���taל!1S\1���9}م.8&�(���gQہJu�"4�l�'��-yW�GHt����[�`�j�����j?��yɭa^��KA>JPK[��]�����'� Dvr�.e�2�TC'�s��?8�ݫ>���Siϱ_{�.�D'x��H�bڎ���J!&�54���KF�q�aO3
D��Y�}���� I�\�\���WY�ks�F�X�Y�?/��.�E�:���ʊ �ZK�^���Y�����v����ݺI�"��ɔ5�cI���}�oND�(��x�jO4��8Y��Cj6}�F�C~�Tz���ikSe�lƞ�:J�	H8��	��#��ϲ��{Y�a�_�[�c�.��h��q�|b��1��̺��%�3I�E�]=���wLESC��U=����i����,��U���нV�Z+��K������9�p3������U6�F\��[/J�[~K bIaF�H�*��ת�qp�9��J�R]p���W�.U׫�R���ٶ<g(y���� �9@����PS_�DJ�����[�I{�KY-��=�,�~D����c�o���Ә0�q+�_�7X	p�����������TX���(dqN2�h,(�A��]���)��|�{�Q�U�I6,���6P�77��#��c���n��O����T7�d�,0C�i`zg��k��Y�8�[�jF��Qf���L�,e.s�ŉ��T�q-W�Na���@�S�!#��u��a��=��w�`�����Se�h��(?�6S��X���e&�V��}�j5b��6�����0�	���J��Ft�@�4��֊{|��>�̟i�� d��9)�����+�kX~i��o�ކdd�}�c v�T��M�A1#^bV8?�5N[ng��j�Ú�?2����8�W�����c���i�gq����~�Ld��"�l;UK�P5LX��:>�*�T�L8�^4r<E0X�b��gw�Zd�^��z��?��8ތ&�_`�Q�ndလ���-��РX⒡�h���5Lj��M	g��Y2�бC1K���*�E�s�f|�	��nϼ��X�ʘ� ʀ����{�cWD�Dh9{ D���}T��f�E��[]5�t"��������]ESЭ�B�<�ch�� U�w����|�HC8e�E���H�a��ʀ�S��r�+C4�w�@����ɪ���[tl�����jmFW�OmeZ��ӱ����#��=M��F߫���b`_Q��v�'�`�q���Qf9���>��(���;��J�Ӊ�Z�ͫ��x-j6��iN-�t�1��	"UN��G�Qv��5���bS�rSjs�+{���Y|���hZg�Y�����=�;Ohђ�J�X�j� ���mM1F��R'٤�n��=(�]�i6m͢�ط��M���B���pF���Ll3i�=��'gX6�.΁{�[�����D���i�(�L9B�c��2x\)�.f�e�{}��>�������)�SC���w�|�Iy�F�%2Ξ�J+��FJ�k��x��x'�E�#���x����Ir<������+�D����ty<F��)XB	�j}/@���8�!��'fl�2��C �qZ��>h�߿��jFh�y"ε��!�떨Sb����љK��OS�gPr*��%3�'zf&0�'[�c�ܦ���<�'��U��	՝����U�Yڋh������g�C���T�V1;�	_�����^�B��-0S���n��׎*o�T��@�(���}Ք�����z|@=S#���`���5I�s�č��9c��O�/gi���;in���d�c���m������z폕����E�֏4G�\}x�5���&�U��R�S7�R퍖��2�'=��j�T����O��p�3�N�����p�|�h$�a�v�P,.TO��T��j	M!��%le�:��؄|�̝��
�pr��;{���1!ҀQ)�Â���03�6��i���¨�����Fl��/�ec`*	_	7���j`�f�u���
j�������_)�6�C�VO�c�F
���N��b��<�/):/A=[&y[O��P&K�my�[�J�W���M����ӌ��{ ���d-�J�Xe*��FX���&���*���C����N.3��"kQ�t��/��p�B�49�u��?��κ`��*�2CR��aE�|{$�dUIu�7r��DS������$X[��32E �=w� �,D�����6ލ��m"�)%���\�n�5�բ`�~.Dr�?�5���_B�z�I�W~�j�@|�UT���3����mh��/_ȳ�����F_`mYJ0��m��pY�٪�2W�g.�����?��ާ���j+�O(D �e�%��,dHz��Y�(T6�������y�k����ޠJ&u��^C*:Vp�Ƿ��״1D_�v�6�������`m��zˀ��QW,����sp���_1��A�Kk����LE�K���z�ɾ�@��ϙjZ2*��cs�8�Her-�@"~�x�7&��$��^�j�&� �F����f�c�=Îƒ���ץx0=���v�a�#����Ue�g?+�7,v]m�k�I����ݬs?0M�}�>�o`ī��9/�|<�e�w5����=��0o�� n�b'����	�����eH�a�Uo1"?��B���!ѐ`⎹��U�̰n<k3ʹ��)��!ʜ5�^m=o�Y��lϬ�V���ƗTϔ�R�QAP��8�x�hQ�2�)�c��N�ȶ�$Eض+k�g�{:&-I\����vo��לJ��|M��� �9����wBW}�c{<��u+&V0ɮ1�NUW�)f��BH�n��0��]/?�^�$��\�g"2����{i9u��)�n���S*IXuc�er�Muߍ�-�Χ���r�:Ӓ!��4ے�n{5�,��O?=IJQ�8��t��x�<Ha;=�{f�Z�H}�[d���<�r�r.���6r;��.��N/J�8�3<��#���t�Ѧ*�>�|��Ɯy���E��֪Į��f�`2Kn���Xf����"�[�*�q���D���pN԰MB�Fh'��$m��xS�-�^BH��rn��앝��m�%�7�� )D�	��.���Q� �w��^���nAm�p���M2��Q�l�4��.P+���Ac�}e�=���[����c�)k�W�沀�~��"]�����G����`s��0,�jY�Ck���/���A�=���E6�vA��5e�� ����:���N��x��ʄ$c�,3�1���_�3��"��B�/:�Hr<!qY>�����J᭡/$��	�X�5&v6^'�=Y�g$����ෛ�6X���������L���`ۭ&\��Q���n3G�TP�BNE��e���<�6ZA�������y:�#�	�����W;C"�cT ���N*FDrlxi����6��!`�yT�w�%�p�X�aQ(U J�w��ߑ���!3�XF���H�mM"�ߣ��M�8#�%w�CH��_1s�9�;/.w��R��Ȯ���{Q��H|FI���⮾ۣgD/�8'�N��3�SF��+z�x?v7� o����No���@��K��.{~��!��@��%���;�C��	
0V��W����2�D{����{��z��]����}+J�b�<�z��~�܏�J�3��Ķ2 ��������B� }d�\W��װ	���Un/�H)x�ŕ�^K���=W�+f{��(����2�L�f1�>��"l\*����W�逴��B{X�/��4#`��I@�jz8��ys��.�E*1�u�t^�ܣ����F�U ��?�������+���:�%[�?�� ��
*�;IA=}�G���A0�J��z��H�O%�3l���c(t|��uޮ��MV2�A��τ�Dqƕ�����jy���e��.����Nt����x �U�^*M	ĮeE�V�!���^y5E���ix�U��5n"�=3Ⱦ$C���g�֐��iJ�����u��3<�������M����=nX5��$|���h�%���7Т���e�a���|���EP�6Q�z&���1��q�y�k\���T�b���(V�'|��ٿ�4@]��t���y������aC@�=w\Q�@����m����q� �:��!֡wx/]ր�nx�̋�i�@���s�Y��1 ���y�x5j������z�`�G+%,C�?���kr�L'����U�J���O�`Pf��7��6.�ѥ=s�����2��m�U~ѵ��W�u�X��g���������<���EK�H�譓��h������2������.,���7U�zMZ'C?X��v�hؐ.2���O��w��D:�3���p�ȳ�p��ȧ����
3Yw���AX<���N���q�~��p�!d|� �k:�a�1�?7j�9.�8�Z�5}E���n�@�u�VOx�Mˉ�F��-�� p���Gm�h��u*��)ʒk􅆕9���q��EOĔ�
&�8��}_T+��]2���D�P�`�\��5DЭW�gIT��,���m&��Ȝ[��v�7����T�o^<{L��� �T1��J��%6�ʽ�rw�y.qE�a����K1���쑝��PE�OOp��V�!�*o�i����v�b5�����"�O'�9Κi�w�9�{�4Lr��9;��t:%B'��ŋc�e'���k�RRC֭fT���~2#�� ���X?�%S\x*�;��9�O��.�Qu�}bmf�������t���ߴ��?7&W�\�kԯ����`%k�T����3��F$���ObI��W0ANSE��?Mbd�-��E]��>e��	x�\6��S�bU�g<�mֲ�J������N�P�W^^M5��9G��s�A��dE��e�D�cl�;�Ǚz7��+�;��<��>�_8�4��
�>*���5w��k��S��ǍvGry(י&����am����X$|˝27��q �y�L��턁�w����-I��Ĥh�![�f��OY�3�ٯC_�=�)��� Y�K-^
�Uc.�h�o�� �\|8�i���5=Yp��D�;P�N)X#����6Z*��\w|(/7���J�Bx���	�w��^=�W�V�m+�\�b�?��q	$U�F~�RD����N�� 0q`*m�IG��b.��O"�A?Q1N��re-�-|�vJ���sK_�у��ke�6�~j�9���[��[�;?��t���4��c�#CP���x�z���.h��:�atb ���xfa���h��LM�
?�#d�oaH��|%l��c��܏K�|��O1��~2�E�k's������d3�8��ͻ������!� Jby-gj�H��S|k�� �e�H�>�U�\2��D )-�Fzt��e}14:�Q�}B1�QГwF��F5汒#r�������$6X*��q�d��3<��ݶC�KaB���h��mr�[�*?�5��@P4���zZ\*Һ�a�q�ϛ����\�EQH�����k���`=qڜ����r��}� �g�K�6�jQ��v	�h�扡�ѓ�W�0㋦�������-ӓS7�b+]E�thF�����O��l����� ��k~O��
R���kY΁���h�m"[,��uqs�ѨHv���jCbrlv���g=R	R��5x�%l�/wҌW����H�5�0�A���9�Ë����E��פEt�&Q�.�2iQy顙Z�Pn�{)��c1:m���l�/�b���'q���1g ȇ�W�M�����e_�1��b^&Nj/�e��3���$aL�������c��E�Q�_��^ϴ�g�F�5�XԮr�7&�֭��%��4A���D@,@�x�>[�`�epe,~E6��p�3�Iv���K�1��H~{zQm�0�7[-P��]'w&#@� e?@������}~��7�����8R�mC�v��	�H��<����]\,v�����y�X�G�,��m��{��:�~Y
R�F��4שf���Z�k�����������%Te�Ϊ�Q�� �m�L!	��2H pu� ������i�r%6Z����m���������hRJ��Y����/M�|�ʓ�9��Y��8-�}���q��I�c�+Z:
1�39�U0*\�c{�)�G:�釟Z�!8�y"@�9
c���v�n�P�6��@�*�O�'�B�ٶ�"���0f����b�����W����	��y�bl������Z�����є���j���>ǩA_#��U*A�O�W��q���]+�쨞if�k�չTE���%���$�#��)�g��t&��/�F7�im�o��y����c���9]I��d����r�N�N�m3XKP����J�֐n��� � `�x�OBj=��N�kϽG�0}U����ٝuIY�z)jמ@ޏ�V��mi����a'�#�BB$r��~S�6�H

A�$�����4����s�J�c�_yrh��ࡔIh�9W�,|�><W��j	�U�ZxQ �^&'?	 �q�n0`��.�<շ�DD�Z���.:�i%w#ʽ����_��j��|�?���O}s݀X�H��G,E<��G���VW�pl=*�\�@�2�K	OM��b�&�*~�'Dw1�g.���[�Q�2O
�Ώ�˅��,�����s��wb�(��}�/��Ɵ��;m`V�>�6`��j�=n^�;�,����콟<2��JU���#�.�:��-.x��_�:x6���RT@�T�>ME?�fe����>aN�j��fQҾ�\T��PxK��{ ?��<0t���'XBLB����4Iw���M�SLO����.��^�@��5�l��Vnw!�����h\tc��~T ��9<	�kr����p����vْA���Ґ�$ƍ�7�J�H_�,�|������t>S�^_v2֭�O��ʚ�M�d%��t�U�\v�9�
��X�ѷ+4
/px�0���9�{�P����*z׊Y�Fݐ���.���[)������$��4�٢�:��I5_L���W��s�r�#�
0�U5�/���D"���R��	���A)������mq���l4ݡSO���y�9�T7CYk�r�c5��`ai��8磐`�,6���	i�[^���n�&�=��'�6�9n�g��<��u<��gu��զL��e~�]y��I��S N��Ť���#ӭz�@PF��C�����eqKC����3��	:�#*:E@_����D#�8U:Фyf��.d�)i��nI��0OC�l�v �bd���3������ˑ��H�O�G�J�9D�-f���+6��<��12�u�)��H��)�UY�۞G[ JD�H�Xx	m���[����q�P�և�ມ�ŒY�;t�ޭz݈�q9D����ѣ����i%�/[��4i���_^M�cr~�Jx܃q�\�g5�"����� ��"���1�y8�K�4�����2�ɮ�/|<Ҏ�>�S̗ӽ����T��]~*VR���� ���$�_i�s��b��A
��:��(�KB+x�S%j] ��u[ɞ���>�g(
'�q�J�ILV䰑��H�Q�'I�n�W�v) ��7~A�P:Լ��|59��7t��L4��B�����i��JC� m�V>�[���S��e�oʻ!��=|'�qб_����o[
�^����C �.Q��à��<2���vy5�=��@����}Z#�D����Y�X��G���/�|
/{&�`yK�j��b�$e��ˋ�ש��HH����)���Q���%|nM��.���!m�5�¸�{�@X F��-��*���=�s���'����Ǹo�h-�+G��(���Hd���B[�BӕCm�3���HJnf0Mf�sE����E�B-T9$���I�S�J��=j���6-�ZC�Eq2��E������vˇv��ܐ4=�Ǭ;�)ә��gg]�Ct������sw��9^+[eHz	���;¼��@��i����Ŕ��c���K���Ϧ�����Z��R|ZKq۷Fu�?EC��=��~�8��O���G����#/�@�G�#��F%���0>��̝d�H�T�U�{�0�n�]����G�i4��H'�4O�T���ދ���4��O	�rF�nT�R�D������̩�rb_5|+=�"s�̵Ol���;�M����˙�]�|N��bƲ�Һ��?r �?��=)m�*����u�P�;���xRW)��_�]'��re���mQ�D�{���j�Z5����Ͽ�C,�~���zȚ��>8�]*�;�f�����%���c��&T��nS�9�.DGA��9L[�}nCnZ��AsI�\S�C���m��M{*9��|.�W��]63?$�k����--�=�v�NH�XC}���[	_�>���˲���}�d�V_�u�����u�ؽ�S6�����,%�evpǩ�hBy�<���rc��l�ڔD#nɉK�a�]0�M��3�#�	Y�ݠU��B�"k}�l���"�4?ٴ=td�8 ����@�+��*O4��l+�^�މʣ.���xNtd���n�X���չ6�9�<�DfEQ^o�ϊo%˘N`2�᪀���d�5���x��$�b֍u˫��Y��y�!5�LGe�Z$~bӻz����:�v�^~%��[��G^#����/��#��*���k�7O\7��ˆ=�=Y�]EG箂���;�c�a�>;�SX`�K��iF:?�	�F'��� <��XK��Zd�/��{�>*c��ɲ,#`,BK�Q����
t8�� 7#�|�Q�U&Ǫ��j�	�b�/�5�/���Նp�#�L:�j�M����|�`�J���4����������+�s5��;8�C[B�*��qJ.+
�\���Nƾ^����x֩K�?�朾�/@�E���R�C�����K��c��QW�1�%G�-��צ�G�U���n���"3�C�{qzO٤�*C�� �Ye_�#*k�v����o�i�m3�:G�u)Z�O��5�$;G}�Ը���q���g�F��k�Î'�0[�� T��$�>l�����g(\�(/y�Q��ohv ��&Wz�=uJX[�<І��p�`���@Z�r�,�|٩���Jw��cZ����� C��GT/��c|婮����ڀ�na��"��,��l²�Z�����nuw�dA:�4ڕ�e�BK<=ӿ?r�����R���#osԋt^(��n�X��{���u��j�.^�Io�?��M�5ɀ� �}}��C��/���?;�J]s._�@k�3�����#ZV��͏��wF�ح�j�V�*4r���.��C��g��ܶ��{�'g�  �����ٻF��z�?�<lTSV4t5i맊SA�Q�$�L�\���Kw�)�hg�i����ؑa�YT_�K��Rr�]��zr3s>�+���Q��].�����|�7�|�̨�����pl{��ΚE-xʲ�{踛'Uw+��4��Pj�u�7>TrE���@�no�p-/�|��u��nA���JQlZ��6��W�B�e�.����H<t#da,�c*r��4�b��c�<� ���ӓ]�<܋����&������wnh�����ԙ"��kI-r+���	�C���W�c�����C�u��]��Qʇ�m��L��ۃ�%3%ƂԘ���<8{>�p���'a���joB�ҽ\�Rn2�<a�U���W8+�I�I�py�����]fo$ϣh�K��#��0oW��}|ȓ���G���P�k�q&�}���2T�za ګK��'R��V9����VE�����Tm:��3�_���a����!�H��u,�_�ϯ8�FI�H��x9�q鵼7�`r�}iպ�[h�J�\�X��_7̨z.%IX�����s#�׼"LՈ�qcsA���z�쟿�`_H����Kyy�����gƛx��)=K��R����V���w�IpI�{]�[l�L��Y�f�ؙ��p@�}0�Wng�1F�~�clzxdθ����S��7X��8Ϗ�X/q9��騖��5���l5�;05nK�?�G3�y�6�0��5���SW�ikc��M,���W��+W��芒�a��Q̔~����/�#r�N�q(���Ww����C���g�k$��`��}��^�_4{���ړ��?G���r��ui��}z��Ŷ�3�F�5�z�\؊f�� ,�>��b��j���37���S4%<M�0�(�pO���&�25=��)��o	����_.�=���7P��T�\8�h�,��Q��Ō�?�9՗���)��d|�d�3���j�5a~�&Ǐ�PދѲ�Q[� �F	[3�CUd��T�t��k��8��E���gI[���r0Ω���|
�lU�� ���yU!5�Z��_�{*'v8�f�x(= �X78�D^�'C��|�>Q�kM�p4�5����� �zx/��awڻ?և��4�3��Eđr��p��o��f��
/���K��IyL��"��.�����LC�����B�ƈ���I��{Q��k�`���D�l ^�C^�6� ���aq�(9��Q�o��!�� RݒDjRm7�c���p��J�rq�I����W
q�V�iXz�b��]��� a�(���+Flb�R�q�yc������s7_T�2M���&Z�tjl2V,������\C�����O��O��E@rbJ!{I�+�g/���ĞIh�,�#��h�+�<�BL
V�I˲̢��-�����b(Øb��l��B��W7;''`$2rR}�ya�������XB��;����B�����(���&�WmسR��9���n����cGR�z�<'ץ-�S�|����T�m�2�;8��f-���=�2�}��{4O����t׊ֆ+ª�FI)D}F��@�쭉�I�Ǌ�^C��|�q�ؾ�Io�d�5C�Q���!� O�	�}�^�ȟw�R��O��	*�ly��@�=����_�̄%�hָ�]��@H�m�`�IW����A��3h�������Ҹ"���H�8�ơ����W�ka��^��0�C݇�lҒ;
�"�=e��<"�7�]� UܹJ�����a���?���:��Tu$�rvg���pR����m5�w/n渋��!V�Tܶ�U��=̍�I���P�胼���"��:ɉ>�(�Rk|�Se���	� �� �R���	,/�>��!Gg��=�NP&��Z�t � <#!��G�q�!S�������ˉ��^�yw=c�8�z]�x��)��Fj���_c[e=�$L��(�:�T���So���ݹ9[MW5��40��M7�}ł'���:cƦңuXӵ�b��,���oBLE_��ϰ�eo��-�7�"@��#�t�,Lw �`�o�l�(�l�o�h�e�ҕCuG����b�J����i�f(%@�N�L�3,!�f6���G�W�/���K �a2��1*��pk��>L�ޘ���͆�d�
��R�3T=��o��'l���m/Jcf6=xz����o�cL��X������@��a]�>2о��^��V�\Jn����tm�h
"z��G������>�:�����Oe��������޶�q��P��J)�8o�S�X$��ar:WE�Y|bT��j�G��đ��\�&zړU$��|g;Z�@�'�J(]-�/�蟩�ޑ��?��S�c�树�2�x��r/���	.3]p�%Ũ<$��s��̑�V�pq5
`<�a�\
='蠏�W$k��ɸ!�Q�:O߼��N��� ղ3^���H�5�[i4P@�Y�o}��$ `9y���t��Y0� (Ϝ:c�L)B9Z�0�&�Q�9��M���t 5Z�$JrF���d�n�N*��ܤ��"7�[�ϖ�ۗ:i�-rtz3���bW���)�@;)�⟂K�O�eM�P�,�
9����I  ��$�Z$a3��uTK�˒�ɉ^}?~vp��,���*$k�tq��I�]�����'�<�=��K�-M�?)�*O��_�x��+�@y��s�+��?�ȁ�!I�g1�"��
<�0z������&c�k�'�ѧ���n��OsJ�&�؝�H����|�.ַv��<uEԥs�{+����㤿���ld�񖈳#�2�!O-��Y��{�O�3y�\��w�/���߂j	��c����så� �a�K��o�� tu�]`��W5�ߏ�G> �$I��4�����}���^���fG�4��U�����-?����;T�?��qQ��'��yzX����Y�!�o[أiN(\���댼V��g�b�1�6���2>��X�b�#�G�RF�3�#bЄl���Ű$���߆4(H��s�3_'��쮁�
|���ʰ����L��PH�f��J���.B:�7�]9 ´3��B��s���� �����M��Jۯ�GF��\3g�ם�*�M��#�ډЄ�V��������=�� �:d?��W��<̛)3us'�q��9��/R�$��[uU	w��kfz�s�ޭ����9���w�&S�^/��|ˤG���$`�>'�c�փ����d�ܺ��`�/�x��+�ĥ\�af�$G(�i)�pmD �ޑ��2.��D��w�R��f�v��x;~^��N��ՎT�`�-o~� ]��Ix�{��[�N��U�X	���q�FM�����ʦV�<s E%R@6g'�*D!��5&q��>�(o��wZ�{���z*��(,5��6{�)��tHK�_+^����zº	3�(c�8��v����~�&�݁��yN@��y��Ψ�c��r��^*/V���'�0�d!P/�*
�݆�Gp�
ޗR�z��x0�k]Q2i�嘎���г�p���jN�f��#�c������4�1��xxŖ���Ŝ�5fv3i����`;�9OtV��#|��D�A�� +r�O\�J8#`��Q���Jł'T���-���\����aN��G��3�ا��#R4F��R`�?�.��v"�@��2F"��E��KY�?36�re[��<��a��^�?aP2��&�����?�^ޅ�����'[�MYм�����'��?�=r�_7贄"�e��ɖ������i̗X��0��=����dY�Sѯs�qڏ�w���L`�E�S)l[�bJ��M�D�Aؑ�=b2���(���)H����^��ӛ�<�i�E/��Ȅ�� ���a��-lM.$c�LE�%�s-�>��ީ
���J�Z['�/�e��M��Ƴ�K���XlX�/�ڵ�w�xf�5�D��_�} !�^�?Y��Hm�B4:\�YQ7y?<�ǈd��WB��i���c�,�i#)j��٨����c��M
>�_ć���=��:��F�=Rf6|?��X�w�4P�4��N���V4�_Bh���o��ٮ#���9lb(�Lm�V�SxV�|\��5A
߄�o���fh�竉��0��2�]��Ǥ~����Y������;�1��.�sv񸻮j�r��8�]�N��KÌj �T4u����`�⸕|'�eW,r^}�u�U�����-]�b>���3��}��BRF�G�f�	9o��~�ߌ�@ �`��+$���s�~h�ad��A�YG�\�R�%c���@�}g�U�k�V�d ��	,�<)�z��FeSn?
d mED&�$��Wk!�s6�ϳc&`.Y�L|ړ"�=z��W�	�A	g���W��	4
��7`\�w���X��/p��3[�7�\���;8��2\�Ǔ�,p��s�]W�n�*z{��zM-g�&|;������!��Ci��(e1��6�<����e���gxEwRS|�o��e�d���������������C�.���EIƧ�=�"](G�s�܎X���<�&�;��@�[�<�$o��f� ��R8����[P�$sl����j�Q�SD/�j�bt�$�_Iu�b8����]ynº�
i�`��ky�4�:?�2,-�Y�G��t�M0k�c���(�q*1��9{P�:�_�Di���⺟."�ۑӮ"��1�K� i��6� �o���y�5��FI ��zDr19g�"�p��t�P�u0I�:y�y�Bc;�'e����WT� \xw%U�{[M�nL�}d���A>N�<�r�	�c!�h��s
|luc�o�A9"l� �?P ��bjn�kN�����y(ͻF/�QBkh�>�5C��J��r�y�E~�U�ղG����������]�8���l��g�)�G�+I�Dr�=B�#uK�jP��)��'iZ�����s��( ��>����TT8=��y�����B	;�LpA'R�'���l�G��a
B� �(�C��Xq���gH�U�V�&@���睚�E���Y�C���B!�g��
�c;k�"��H��9�:`)x񄢡k�Z�qV��^#�zeq
�M^�h��`W��i����ϢJ9�2O�cfvˊ�fA�.�g�P~oT��X�)^/���dN�i�F�ˏ��2._�є�68@ȥ{�X�m�"�<aE�@��O?rS��B� ݜ��3?g�xI����݋���,P�d`VS���W����\F�^/G�oB�֥���X+�xU�K#>
�RP�Sv��?����▱"��G��/��j�����S�*{��I�!V�~����D���C]��ܹH��p�4I~9b�;7���(�hz�� *��>u�Z
Z�I��.�|���%��hv�vZU �|0\��UL7qj
T� �b�cy�%iɮ���zQJ+��X�.�O"��L�'����g�K�T��7;F�(�� ���F��x��W+�h��޹���z����lbtj�OƬ�B���s�t1������=�E�Mš��M��V7�-�
k�K��^�>bX;lX�EX5�#�`��,��$\:f���kny�t�p��1N���a��][��5��~�񏥔�"��Mť<^��}8&УW��z�L���䄫�k&�?iG�K�%ˑ���]��d��0��Pǚ�|=�&��͔vL��'�� �"02tE�/��c�w E<Z�@�x3�Vsp�])!i��L֠��ejx�,�'q	e�������@��҃ �9�d����j��6��=X��n察lGd:2"��Bb*>��r�A4�ܰ�)�A>����`�#]�j�����V�����:��ǧ���~;[J(D0�ԇ�J�~�Gk恩1�X���be:�kNJ��s����;g�h���哼��<l��o���J�E�vF�kBx�� c�HvT���q�M�w�=�cN��8a����A�
��j�HM��\Y��M��a�C��� �L�[�}vj��|UQ̲k����l�L�Q�r�-��P�頄�w	��fF�ڏ�y��ǜ��T�(3my�'+��O�O����;b�t�Ϻ7o�D+�u��`v��'!�E�p���J�q'��F=��H�f�h�GZ�ר���X%⑵R H�T���t%r�G5�3���Ʊ�`��������jU�*p�P9�3(�{ �VWw�u�u�
O �үT�qe�l�r�'�M��6��܎�b��4j�нv��)�l�^a�0�h�k@�@��W�*	%��}��׼�sT:�Rn{�sdЎь��c����dC}�q�]|�qڍl���ﭿ!�܍%CT�ɸn�
�_�֌)!%�~�{ϩ�E}�
9\ �B�/Q�<����&�:���:��ޟ�������w��&Fb��,+� ���5��KQ���,R�t�=$�&n��+�8-����7���9��cz;����'��h�;�2>E"ʙ�c϶4v0���0����;�,ᘝQ*^��I��-Br3�3���DM=�Ƭ5�.c�ܖd��j�f�����rOL�{1�E��\���<@e�$	)�N_����jQ�&����C���XIK�W���7�fp�!d�b�*�������X�[�����b��0	ۍ:���j6]�8��r��e�f�[��}��x�B��,����f�\f�L<gž7��N����[6� Ze\�?���'����ʚ�F���;g�E2�8Q�������kɎ�]�̈́�W BMk2՛Y�
��s��y>�j�Xi�ټ�S���]�Fa�K�̅�n0�6�J����:>�ʞ�����+��d�a�ͭ�ʠ������ ̼�I���7%�-�@�3cN���K��<P�g�����=.i�+��bd��L䦪�~��;_�~Њ ִf�j��&�s�lٷ�pd=`<�2_�p���u���/"����FYu+0&��\�|(14�lY�GJ1� \��h��Ĵ����l[�"<�` UϤ��H��y�*)���k�&Q�J`ͱM�WC��ͮYy�������zV��͠�:" _�z��lձ�=&������m�Ԍu�Jy,�ץ�F%|��F���1�Vw�}�� ~̢K�,��4Gp�&Sk�����*�&��.���5�����mg��Ky�>C�o���!�����0�J1]�U{\�D�N�$��#w �b�+�����pH�"�5iC�S����yh�������͂V��ƥ!�+���@<�"#w@��$����~�i�4q�G�P	���إ/̂���o���%��A/n�8�4!��%2\��	��I���ү��Wf�p�1h����L	9�S�f@Bk?z�g���E[�s4Qq��loz����M�z�t	�]P�x������(:q��>��7����d�^ �N�E�U%��ٰ	�Ȗ���OŔm�;d�Q��E#��+��U��*R�� �(slH_��<���,�ɎBD�H^ܮv���oÊ�_m\M��/� ���j��߶��M,�+���X���?���W�u��E�#��:'��c��"HOd�r�2���0ش�|�mc̶���1���S�A)/�Ɗek�(=�nJ�Yggh��]�������0s-[�%�g7�+d��%�I��*�����v�9ཊ�h��E�P�^��{�s'�挭,��@4� s�qF4�6B(���ֶ��u�ti�)��
�p/0g�i�[�A�\g�/B�[U:*P�m@m!Gp�Ɛ�_����=�I���?�-��&+����2�r��ף.���ƞ��|�l[B��eȪ���S��hc�Nqӳ��N?J�b��i�qcg���Y��1L������>C&��4�ۧ	��u*Y��V�	ʉq>c�~ה���ba�� q
_�X�-�Ã-�Jߖ؂�*i6��͝�$԰�������KI����X�EG̘;C�B���ȏaQ�[12����VSޝ�+̣�.E����.�����H	b0�����5�O*�(cH��w'��������y�2&����Y� ���	��q�8�18W�˙�-��JA޳�NR�p#����q�8켔i�"x`�Gh�M B�~���恲ˠ�2��΅/;�1��(сS'h7�n��}}NM���R���{P�a����Ob�f���Ҟ�x��u�Axz�	����2;�&�E���`�ą5W��ѳG��Y��� 6����rk�tЄl2�O5睇��lU���@������v�\�e�ҥ,��Co��hZ-P�KR������,�N<f��4�V�'���&vT�����	������)j���_���S��~�T�q4.A�m���*.Om��C�����l�ݏ;�8�v��b��ռ��\�!�������-��"�ǠEl�W��{���Pj=Q�qA�;_�UI��?�&�nq#1NkL�QSѵ�����k%��:PnƑ����٭>��X���kx��l��ə3�^�s6}�R㥮��~���a�/�>b^�>i���,��bc8y ӵ�lyи[�h��kv�큋W��I�*բ�0[z�>I�}q�c�'��1R'Q�����m��U���D{!�{�cG���;Lx>k�f*1~VFi�v/��Z��ċ]�3���KS r���!v����=S:!N��<�`u&���Z���Y��W���Q���m�[��l��J��b��s�ב�Ot�����
���}HMSm����&�*��ln�=�1Ź���.�_7����Nc��s�`����������1�XµP%�9M�ه�=х�_�h��Tp�
Bd}:��.��B0��u�e��䄋K&�f/�/#��D��8�������3)\��3�29��>Tn��V`���D ������t��}��v�5�gh%��O�p�+�I����la�T|�8j��x�tGM���2H�z�ſ����E�?H���'��#����̪���ì�z���N��!���Ǫ�&��"���c�=ED:$�̇�E�@��%�K*EwKp�b4�4�Jv��N��â��A�c�l|�f>���,IY]��x�	����{��?˰��>����Zzۯ@�YvG9�\�d�_���#X��,D�"V�����yX�WxDЙp���'8{���n�������O%�.�H��!m�R�fnM�τt�%kD�ܜS������7�+�}O�D���J�o]Oa��k*r���~T�G
>�Am�u��a��U���tP��IE���Ǽ_�6,�7��EO���yw������~�@<�F��'=Xo)�o6g��!E���T��T4���dJq�5��q���֡��.��\�T��G����,~�s���k��e�Y?�4�9�*exG������n�-|!"	��}�+���SA���r��:Hܹ� �As�KY�8)QI�2�j���rY�0R�$�Y���s	H%?��NV�N䚪��)7�#�9W�4��["�*{��.T�18A��|
W�-h,Q�ԓץ�Wel���WDp�6��s�0�.�����J�~r����C��}�+����a,�U��P�0��o���Ê�!�����#������1����v�5nN�쒞��%�yz��Ř����%:aB�?P��gTk)�6~��]VЈ�1۫�
��O�+��hӹKd_�*�T�RF��A	��r�xu\��~O� ��l2̮�p�~��Un�d39��)�[<�����k{1�c�JM�x19�鸉=�6v����[���ָdv���w�5�Y�E���:��h���4��O���b��.�1[��+���������]���Qk��Sd��},�;���H�/��h�F�oC1<5=uF$���$p;Y?� �iR̼�
9^��вʽ1�Mm_[������נ�_m3��x�Tp]�i��]�_ �}����@yzQn��f����J�M��A��L��-"�g�Z���<�M̜_1���C"}��TQ�6 )�!dʃ�3��#_-���!&���ط}t;��S@(�|P�v���L�7����(���T���Ñx_�W�����=�P��5����y+Xw|�7+\�n��'���,Ql���;"��D'����VGQ=���E��A�L��M�����/:&_9	��J_y�� :��+t?8��i���~�#��Ux_%X����e���zA �J.0(?H1��&�w�����K�Ϗ��+&��cP��Z�@;b�e`�ㄈkl	��c����[7%�d�k�%>�TD\�}<���5�c�8լ����w{g����R�����o/� Rp���<�D�k��I�hSL��}�u K�y`�198�������ғkЇ�<�B��xo�����-�:g˳�^��W˥0���89�_V��}�;���M���gW��n_�L?O��Qۙ�.��/n������5�}-��F�iT�C��&�o;>�Uh�H2�M��a���f+�-#��u��'[�2��z?���҇M9n��i�
�M�/������Ny��6�%��L9Bb����9������`�|�wr��+L��W���u�oiP��ʖ�`�������>K�J1ү�o��E��g�*�cK�.��
RTr��fĝ&Ȳ��5'�p�$�:2TBr$O��F(ʺ���Ox���	��6L��/�Z��KZ��E&� `*#�"��%I�wM]���2l��r� Cl�|��ۧ����me�l�
z+����'�C��En��#�;y�{Hj�up`�YV/����˘F<N�H��7T�dn=���ܜ��Ǧ�n���gw:�W�*��[݀��1�EI�	�xG�)&�̠>vn�4�==;�7m��8`���X��=ߣ���.��[̂rd�{l
�j`�q3گ�N3e�X�Ժ(�\��
!�{n,wk����9�A�,$��r���c���y��^O�&X��ar�:*�k�	����9^E+����|�ȗ�ނ��G��5���\���_D�Ǔ�e���N�g�m�����q�7ƪB�R�:��^��f\{���-B���(��0BtB�Bc��P�+�oI	p��m�}���!��_�n���'s� ����WY-&�oZ��^�-��T���i0����	��懴��l�3�l,��)3.ӗ!�阖��`���R؋�P2e!�YG��-a^�T�˵� ��"���9ʳI��ab�N�ֶ��A��Q%!��b�I(�F����y����_�]ݢq�֜����N]����g�+a�_L�L��.6���Z�!V-�j���Z�]qa՛p>X�O�,��q��C����W<�����?5��C�x��;⑄�[y�a�Whg����7���е4JK3YP.EΊ�6;�����J�U�x.Q����F���~|L�#��	v"�$zZ`w���n( "]:�Q����<_R���0�Zn�gu��<���\r	�`�p�|�߇����,���ϯ'� ��弌+O���NG���Š���^�u0���f�QT%���I�=5��C�r�_���(�q���s�����un_n�\cA�<@�e�ҙI��V:K,T�����Go��C|섰 ��o��sv����ѡ�s��"em�ݪ�r��*W�!VԳa� �C9���p��3�Y�Y�����cXH���/.�YՀ�0'r�G�4�3~y�HyUc�ΥgK��G#l��G�*s�&�d �t�Ksj>Zê��ʏ�v(DV����bh2]PL�������gp8��oqݹN��6��-rl)�'
+���*����1v�Ыk�A�X�H�)�&���5P���R���ۊ�cR�K'�!���ȣPYxa��'���0�
�����f(��&Ø���VbŦ`G���'q5@��+����K�l�-l�U.�(�����o���裯F�i�F���)Ct�����aD��A�e
�j��?JIT,��
�o\
Ɋ%%�z�}*��b>|hGI��)�{:�'�ԍ�6O[U�O���*�|�s7Ȣ'�	��R�����Z��$��v !p7*����m�]]~e���$LGg]:�C��s�FG�K�0>6@#��d��
�n��&�/��}��ؤ�k���?6<_�[��ED鴟{�M���8��v�^f�ģ�3�r�
���� +��A�}��g,��J�l?�^���l��6B$�ԗJ9�aLM6n�F_�XA����'q�ѯ���p�p��͏��\s�Q��^�|��,��%d&q���]�8�.o�t�ڣ�C�5�ff>������f����_�T�Ք�<pR1�2X�x�$��ů?�τh�,��Jy����w$�N��7��L,X�Q�X��8���ƚG%�G;"!
��#�n��˱�5ڵ�{
�c���5�����/BRK�a<��\������Pv�������_;n�}P�UWmhO��UO���I�SEX��O,K�/���@ˉ>F���2֧s)MTmZ$��q�[��������0F��t���@FG��wu�+w�o��K�i~���]���i���Vޘ�F�����
��Qa}H��$���+x�|��MDH���n��qʛ3�|ΎܗF��+���g^���6r�ja����;�$��<Ԕ�o ,	��!q�8�0��-L��W-v���ٗ�Z�����Dbk4��y�Zt8g{����}��W����E�Px��"�*�NC��Ewe�\�C{$
r(�v5��EDQU/2����*,�z-�ay��|h������?�D/V�s�G�v/��%sk(BO;�
�Tŭ��^�iGr�h6�V	���l�i�,|���n�
�Y#�L5�	��%p�*��&�/���+y�A��|���Hl�"���Y�D~M_�E��=�k&�߸n�]��uNmM���I�:��&�='e[s�����8���^�w��l�X����t=|_3,|�l1��YK�-��⼖u�V�Sa�<���<
�K��T[���/СX��� ���3��ul,A4����x%*�R�6�}=��9�S,m.��&f�ྣV�U!d�-~��jGU��䕨Qt�{�o���{9��(��q>W�׏���<o�����IZ|���N^!��>���C6*qߊWV�d&ҫ�&�?����u�=L�	��iWz�q���@1D�ZvU�V�י���y���������t	ׇ���?��v1���d}>l��$!ũ�2\�4��c��S�ϋ#��=����$(��Z-�xt`�j���-�O��z�f6���~J!H߈l��qr�,�E���,���G,�]�I�T~B5�)Ŗj�"�,J�ޕ��[i�G�!�q>�!^�G�<~!p��o_*b��jZж�EƘ�a&�Tǧ�+e����CGʴq�')�LT���O�	d)�~����0�襷����M*�U��3�vE�S�����o)���,I��`4'�d����W��F�D�;wzA_�� �uBT��UOj���M������|6jQ�3`_�71�&��C���%LH�q>���M-TM#�Y�Z�ۧiJ�&�Og͘�)�u���6��<�7��OL�*�zZe�s����3���T�P�*���͇/��:�=� 8C����jQT��aV1rƎ&Vq�F}"�Ӷ��贀��}��K���ut���pIc�������~9�"^Z��u������h� ?���I��=�� aHZ�����(�����ٚ�U�lzf�t��N�1	�E�F��g�'���mt���R�"{G�Z ���v��4[c��21�!)̈xN�u#�q���asn��GFښA����ք�`��HD�@k�^ͺ#�v~,�}��_�-İ���s_M��_OB���#�\z�����X�O�MnJ!�t�Oww�1@�����%�����y��sk�!�CGX` �DJ_���L*�!]��W3BP�P�\�Va��8�$+PA)~:���^{u̝���,cL>Wm�3aU�����X�p�
[�͑yF��E�	B��`�NޙW'�%*��+���>��
�Qv��9؞$���]2D�<BHg�5�u�E$g��M}w�s�1���X�D��](�������*a��w�g�����i�� ,J��� ��b���_[ Mw�n�����v�є܂�ј(��'Z� 3MW�<h���-_*'���V�W��gZ�g�I���+�P�����V�ºd������E�g?J���R��r_um~F".��?�+M�Q��S���]d����?/��?`�s^�*�G`v=�Gu�R��j�%�{y't-�j�J�Q
�E�>;�#q����Q��Ǥ�l2R��
�K3JVVZ���%e\U�#�<}_�����K�Z��E��ћN4�w�Ü�#���`�̋�sw��@9�s��!F��e vrG��.�=6P KPJ�����ǟ�\(�B������p@��^��^ �d�"���;�*�TE�,�-���������׻����.0?X.��6&��*T�?�|���1��,��[c�H�[��g+�+�l"u�C��:	3���W��>����eNI���JH�B�J%/̨+T��R�����@6��?���ƽC� `����	��D3RA��G~`�Q��<�����4	�C��A��`�-�E�Mq���s�]��^�T?�;�-���^=E	h�i~�C��.��̏�ʪޔ\�m�o�b��^k�{|��aiJ��F�zaמ]����u(����pU<ղ^(ys�)�0z����RQh
�˛��/'/�����v���Yn}˛��������G��tPL���Ƕ���/�`U���@	���vů�&�ٷ� �����S[{g�>,MU0w�`+�]�D��z��*����`��h���e���?�/:��C��q>�G� 1�z��: Q�oN��Vk5�}I�[�)Eo$Mn�?-�7�^�q��kbq�%��a
�g���8!�#�4�5|�2b�>��(:��t�����o�+Ѭ�sC�"Q`�8����r�Z�a${h�(��1D�\�Ǭ�W�A[�Ō�HY��|Fk�j�T���:�6� 	i���ܙ�\$p�k�z�}t����PxNd'����D�#�!��E�#��Ľ���|�:�p���n��m�d|-O,ʇ4E��ϖp	[H+A29�Y���̆!�Da���=����;d�ɟh�{�_�ʘJ{��Y�
������n1e�+d[�㦰�>�x�?�e7`��%	q+{Wj*����7�B<Յ�g�_>-�DgG}cB�Z�ƻ4����4�;���l��\m�<�֨��j"�(����$~���+�z��O��,�ɖ�E�����Y�vh>c�:�����W���Z@��x�6}����z�pt��r\O/
�1����$>%����,�6�Կ��l�N۷�� J��%�t��JM�P1A����c�l��
�J��F�UN��T�)A�.+l��oF���qU��)4z�)ހ�Df���b_��9f�Z2����2��8� 00��(I��O����o^c��G=Cc񆿆��"�]�@�n,�b|�`I�V��Һ����#�����>J���"BY�z;(s�<�e%W�*�_��l!�- �yx��[��cQ���_�l$4�@[����N`�P��;y��Z��%���Km�8
yh��<IѢ�3Y�i>j���Y��f`��Lu�*Q�QL�扆[�g{eU	$h����ڕ$��T�i�R����b�8�>����4y 7V]r���c���Jg�}�Lp��)F��a�_�h�u$��<I56�I�B������o��2��) ����1v�Вg�^;C�O�iO�����=���%���QK�jv;��.�;���ޯ�M�ӣ��|U�t�e@�@���rM��J���z&�N `gu:��E�6�F�ܳ���+��;�5\�/���t�@�0����c�:l{����Q��ܤC&3bI�j�86w�@�����R����:���f�,��=��57Y���j��s{Ԅo�"�GH���q�0L���Q�G֢ap�"۞]�\��=mi$��t����X����=L�T�����9@8!$Ȁ_�)�}�Т��2�R�����9�o�L�w,?H\X���]�Yc8K0#�1�ׅZ�����6 ɣ����d�7S�wPbc�����w�m�+^Փ�0ޭ�p��:���.� 9�Y��!?��0g�.�bc^\�,�b^��3D8�m���/��H~�t��l��ϐ���=pQ����XsXW귀0k�/o���w�g�����D�'�櫥��P�B�Ǿ}1�gF*Xnf��
'���UCSboq��&ox�M0՝��Qj�I�H���2�OH�ڷt�wd��MV�F�<`��=t�,OQ��B�GŮ�B��t`3�	m���(/��S�ӑҺ��Y� �P^Q�ڷP����)W?P���j��~af|�=26c\u<�yA���v���{%�D���Fd��Vrj���!��U���a������!�Ko8��&�쁈1QOT��e ���v�%{ֽ�T�-[T�V�6NhQ�R�����9��t�S�7vbZ핮~NƗ+'bu�A�wJ��F���;F���m��n�Z�>�b�׌3<v�}k�}"�K�G{���K�wZ���Ųi&g���M|��=0�p0Y0*��Ƨ_`�Z�"?t	+�g���'�T��DCd?6Ҭ�-8^�f��M�{�V���I�Ȃ�-�d�~C״V����o����=�%��?�XVY:&���)3��S>a�I�ι3�d��#Zs*a�z��8��tr�!O_�L�r��I`��±>&?I��^��Jv�����T��+��&��8�n�'&�n�{��dj�H����I⬖�M'���Pq ���5H�y��"���^�ӄ�"!r���[��,X�H��;Of��P̲�a�o�aY�ŏ{�a�����`�i���B�RlS�uD���m�}R�,�d<񫴼$�bK����c7�c���,�(:���5�ä�Ox��VPb�RJ"��'��m�-�Ņ�"�6�7�K�{p��r����b��� �j������<�!fvs����'r}q��"{*h�;Rΰ^�v�>ֳ#�F�����pj�Z���z賮�_z:1om��t�=�}�bt��{8�RD�@@�A��by����j�N�gx���G��>ݽ���ڷ�LY�P�� ����B7�,��MmqW���/(���ܔG"�o�'p�{.��L�hlC���-CN˫?�MI�܏|���/�o��g�1�"�yҙ��I�h�ͪ��Ȏ�N�U�U�:��n{r�Y���B����x��Q�m�yJ��w����"�t�:5�2���i��8=K�����������)~^�=��L�0���jJ��G�ӕq��D/��B��`�e�P�[����'eES��T$����1کˣ��O��oTTp����g���D��PB�!r�D�Hݷ�z$d'�m6��%�/n;y�b�z=�.ԂS��P��H�}T�d<��wu���2)HF8���:y��`W�K��W�N�����e��|�]ɥ@K��u�������u"�]�C쥘���ڀ��5��2�"��'U6h.L$+)��k��R�>�����c45Pg0�M���o�o��@ )n�ٖ2Z�Zw�c�9�k[��V�5�ͧ�)mE6".+����(�CW���ζ��ﮍꌀ�b`7�vq"��wM��+��&�\�r�9���t\@�A� ���WA����%?�E~���o6ݘ�
��5�L������@�uŮ�n'8��m6Fh���Ý�PLM؍l˹
Cl���F��}�:�"_;L6����HG�ư0�c%�2ԑ�;��.��,�������=�=LZ��-2,XP�[M���e8%$���G�r�2�A�C��T�D&"�O�r���nz�s���FG�*69Q΅)�`O���g�F$��u�����Xa��|%�aV*M�|�\�	�X�<=��V�R,�ߖa��qjt�����TFF �W�m���զ�":��/�h����5�-{D�����ͪw��F�^y�b�S��U` �/�Nv�J��v���⍴��֌����C+�Ӥ�c��H�@��q�
�Y�bs����4��.#9J�C�^��V��<R5�붔�J�z8e:��r���1G�j�Qh�A�Ҙ��\�:���NOp	�x� �����z�������M��� 7�R��]���@ԛp�iD!�Ļ���RjF�0�/�Q�2��5���6[��2�M��vI'��r�_��4��Q�-N�;��!����V�D/��.&�=��`�M�6��l?�ϡ�na0�4��j۱ՍJ����Iq8�&�6G�B^H�o�+��1�	�6��a���Ϊ�8���Aub���au��C;����>�mZ����M�\��*{�Ԃu��(���ܣ�3z2�`��;=�������J�UF�;�((��w[�fm�GT�����(2��Zz�.8Zp#~��?�*)�?��_9�7ͩ��J��~!����g<*�0'6\SZ��$[��c��L���4|�	�@mW]�G���sL�W��g�ܼ	3�a�N�t�X�.�u:�~��<�m{C� �`�������$X�]*(%wC�0��&(?���H���#���X,�8J*���r#�������+��ȉ��ѫ@ݎE� �>G9]�\��c���S�AJ:�,�n黯����6��2$�<8������ac��qdM�O����O��i'A������~ӛ<N*�[yg+WD�:;k��\Q>�Ԥ<�0��}C���&���/]��EL�NW֕�ڲD���f�hZ��Ʒ�>W�g'оvz��'��S����	_�:����1=x�,�F��WL,7FI�~�fM�K7�w=����mc6P�*�h������v͉�ȝ
�����x��fD��x;�����-P��aY�k����\
�i��:���������v�E��#����*"�04�W�W�9��<�kEd�B�$rC���u�*����Z��|]�i�n9�֤�q�ҭ�/�a�_=�a�D�X�gex���Lf��s�
ըv|P���F~��(P�FX8�(�����j��`x9��n�x�@�z��&Z��ȸ��SYTk��_����ؿI���Z*�O���B�:�љ����̅�L�����.����h�&�r²��$����@[&e#�!SNH�\bC&��2Zy��K!m;zD[�b�x^)D�ӄIuI���>f�2�P��A����ڰkr�0�{�Ȉ(���e���,�5��%�l/�� ��X����Z�G��[l�;:�(�V��f�O"L��؏1s6���A�ĵ������8�^�E�ش�`��%�������#�RZ�������\E{�ݙ��t�z�l$qEI"�o�F�o� ���NrO�0Vv���E��U�(��+׏z�'��/#��iqw'�V?��8 Q�p���f���ÿ��x5��g�;-��L��00����f3��f�����à��W	��Ǆ�j�&=��?=������u�	�j^���s�0�=&�[�
�t]F�Q�Cy�='��q�%��E��|<�4�f0�	����%�A�4�\�p�ڄ0��S~�{X�LY��`9�������\%)�󟤿�A��/Kp]�{qP�Wޝ���U��Tw5��v����^�P���[ŰŨ�oC��!�FaL�@�,�s�z��t���j�� ]�g�=�䭓65�ɇ��|����P�"�P0�af�������5�R��)_#n�:�o�B	��3���|E�:��ET�Z�%�㌹]f0N&�d���![�.�i�8U��6�I�0�,l&���Ҹh�Ka��0�������J}�g�5RG���sS���S%M�@yƲ �9T�L}���b���tֻ<k��l�%�Tl�� b6�(��C+��i<���91	"� |g|J��&Ҳ*6��ji N�fW�@�H	�ƁYD�|AH���6k�;Pp�~�4��� �h[p��*V���۞z���	��s_�+1�{�,j�	��
��ˆQgIb��x��I�RpK2Ʀ�%�)��U�dT�:ݰ&Z���O���^ �[	NV~�Y`��4�u��N׃]��
���XiP���3�;H����X�ԁ-6�C�?B`=��eqV�& ��1o���������tL]\>s�6{�A��sz��UP�G�p�l��s�����2Z�0V�/_9���=����q�Vl�'F#n1��^Dq`������T��@���]ĺ縉.'AW��b��9�W�]Eey�U�h�c�}�M����&�aM��.�*_���2$3��!���	B?;*�:�X�4��F��y@���3n?�t�.�LJ�t������:���fό|XژJ-
����(J�t�q�"�`u�諚�hM�x����<�H6�ʹWR�
t�O�%�b�� �]o~tv޽�H\.���S��Dgyؔ�ym��߶"�o5����l
tC����DP�(j���˓ �� ������zNAJ��π�c�#[W[V����9YJ�����H�=��%����#V�K�@	a��$�+FӽLLmtu����y� �n�o��{�@���*ُ�-�@��ň�k~QpF�m�E�(�J���]W��7����������ş���Y5)d��9)>��������@K^>�\���gU})پ�{?��VbP7a6�nY�y�林��G���F����L	����bu�G�h�[�p-��<�"љc�`S��I�HQ��|�_9ky3�!&��k%0��o�a��nC��������*� ���x]銌�*$�E���^�o��f�hW����kD�J6@򑘠�s�����iF�)Q\�EJ�q�ҏ����6����|gQ�Y�|��{�ê�Y&�v���%ϞQi�����T���fe�D�H�^���	2���b��z�/
_�r�EV�,�e��6�v����`:��q�-�|��2��~�M(P��!�F���+!�թ���P�|I�z���i����>eیj/_S��MɊxE<�@�&e� \�N�㥑C_�"?�E�3^��|���u�۝TB3�J���HN`h&6���MI�&wDgo���sK�H�$Sk�~��4y��O!�Q�9�;��r~�o��v_��m�!�������w:!\M�����w0�l��kw��
�M�M
��MY)��^Җ?��:�,V^�-A���T���w��$���c2�� Y���	��
y���ܦ���q7�r,"���Cau�˶s������
r�҈��ۅ]
~�>�-}drsH+���s�����k��=v��U��	mCg2��=)t|�s9<�'�C�l쑳]�N����wWoS#��L��ŋ�ƴ�qR)���\i�����1�W��,7B6R�9W�ܗ�T,u7�N���6�.
�����]�b��guU���h�3��VE�Cg�0~��_FՃڅQ���ی���HF��Y��Śڵ�Ih8fGƳ:S\�Q�E�vC.e���+�h��P,�E�c<e t�~b����nl�hU/M��@XnV�,�0��vrfcWHp��=������dF�[I����a�[�	_'��'��2vY�8;+~.[
�v|���-��2.�S�K�v��b�vM敀rgs>���g)X02NM~�C�����啧�2
q,�R�:�J&��g����mҳ��Y��<]��2�qU-7�I{��'bI�ff$I�\3��������G���ܒ�ǀ�9��`���=4<�Vŷe9��e�ڂŨlOD�tcl�>{*-���u`+���D�.�i}��+�k���N���F��ߖ��}����Q�ճ�N��8!� �N��?���P�m\4`w�J&�����劮ǰX/��v�F_۬�T'�`�<�أ%�?�����c� %��:^ڨ���9kx��M�����Y�#��M-�Py]�Iܣ(�G�v.\PЄ/��R:~�Z$��r�k-e#Λ����0����%�[���7����/��8Q�\��ZU�AI���4,0a����~Q���wYP�����x��^U1?����_�N�k�<�ﳔ���$��5L��Lo]��d�+M��uI�(;�96���#0~��o�̴�9�7DqS�5q޴.{*�K����( ��:���V�Fɹ��e�����P��"�:s���Y[���6�8�데Vä�W���0���>̭���i�m ����#b�2ː��1�k�Z�c�	/����e�_^Jm���`�τ�<s�U����甄�H#�A�{���!������+���6�+Ӎ0��yjM+١�x	���;r���U���?�W���5P��[dmA���\�z���D�|ȘɛNr�>��+�M�|���
)6mw��8���8*P� �����X��Қ�ɉ��hQ��R���S�M߯�[���v�#���x��:%D���p�L�KIs�x..��@u�e��F�/L;D��7��1&�q������� `?��.˳v�ð���-���_2�l@�:��d��,m7�gOȺ������B��6�8���`�;5$��N���"�V=H�����8��츬�Ii3�����L��!Rw����R��䥩2��73�*��&�Pt��ӡ��r:[�s����u��D�:�A���WL�Ͳ�	6l�r{��}:b/��)�D)�-�X�^j����w�@�'o���u�	����ghX�}�����Z�3� }�XTvc��B�6���=F�!g��;ۧz�
���u/�5�IP���	N�X�[�BDg?>߈�]��	m����m#
]�}-�yI��_ʠs�+���J-t�Wrb�1�b�ȷ�L0��=%�t��Ұ$ď���2 Ҕ����|�C½��R�!1=���e�=���:���-��*o��^�AM	[:�wF&ka}�6gq���MdH��L�����T��%T���>�F��>`�o9u'c�{D����{� ���c��G�Y�Bf�Y�MX��D����laEXۅZ7�D��wK�3�V�$�,�&�0�7��m�K:\M�hT�[��0� ��uJcT���~
�m���Os��C�K�
��&�J��kr��{*���juT/T�dWnT��bx�Ug�c��MoD�2�v�d2y�ޡ"�~��+��������矷�B�\��'5k7��¦��4��<ٴ��"	G����ŀ�+k�tA#V�6�~h68!2ؘ��6ۧ<��$���Z.Z-2����Os��2_������D�ޔы�N���[�_��uSU���jy�I���$�;z�/�j�=��S���z�$R�h��;�{�ƣ��v>��tuS����X��<IoL�q������cBjM�R���?���'��p�v=p5��z�,��L�M��~+X��ï���m����.{:���T/��v4]>ǽ�R6p��RER�F{���%ӭ��=�&�!����K�/��+��n�������>qy�����S�������������/X��6R���5N��QzR�����jGz0���8w��߻0�����e�~�� �h���
�'!���1[�,m� +�)���%!�?U�ʹ}�A�U%.RM�I�CJ[b� ,�����:�	���o�#S����r��B���	�����<\��~��Ӆ�!��	b�b�2��s'�M�9���9�@��/��&L�l�v�!G�)9�8�Ϳ��'����`f��x)��]��G�^�ñe�Ub��p9� QRuΊ������Z!$  2������]p;*�3��L(�&��56⮪�}T���0"���2�^���_�6���K�JVI�g�`yc�[�PNIui���U�m�T��/P�����n�	�-9.�JHK�u)��JIoHC�R�v��#h���<��2P�H�ꦴ=<q��D�		(��e����!Xo&y�PVy�
=jz�@�.Xb��c�m�|k�(e�7@��.��sq'-(�On}�ջG��N�|4����EZ�����8D5a����!�O����o�P�Y�w"�,͎��&6ƪ�7ظNjF|��~7���Lz�6���ɺ
t0:ԛ��XLG�r6Ź�ڢc훚Nr7j���y�0��eK�̌��V�n�����!i���YL�{
�G���<uÞ�u]]$u}i�L�׸����#ez��oh���u������RLTT�m��T��Y�@�W�M@M���Xo�,��o�i�h��;L�{tqkk���
4	w��9XdPU?F5#�S�K�Tt�go��,t�A]��:j�'���R(�X�����N�P{���n0Q͈'L�ă4z�xX,^�5Ζ��9!1!�E61�x�o�j$�}ܐ�����Ak���L�g�$�����S2&�_a%���
���[Q�>��XѠ�<�e� 5� �B��Դ�o�hz���q�M�����o�=���i���(�k�ۂn˜wq[�&H��#x8�j�� �y
~���u�.�S/b���<<p�+7>��,͉��rHz��|���U'M,�T���9=��7�f��ϸ�֩�����ڊ�q	LP0����~5 "m���
�rŃ����D�����8.ߐ�Cs�}�56����z�Av�x�][����\��qH�����(>+)��FonT�q8+0{O���B2��jb�g�Y���ߢ2B|�T�[m�a;�C�=�tBT��h�å��H�M��1��3n�� ��G�'	��4�YĪ%׼tD�I��Ř�6�L����3ߕ�Xy�e9R6�1����gi8G�D��m&S�?T�_)a���"�8���'�]"l_�f	�����-�⟱Zq��	�:C�B=��g^&���@&x�0��Z��3� ��6>=;�,b1+YB��F{�������kז�1�Ja�T;�g��B�4[�q�VT�@�'~��Q�c"�7o~WS
8K���P�Jl�E���s՜߬�|S~r�&�bzD�l��|/���+�HI��=���@���N- �3����h$3�.r7ܚ���?g�z�1ey#��&$��!�����n6;l��ML̷����&�\q�lR�K�VX�M�F�'Wi�`1TEem�A¿M ��wJ33g��G0C�1,�wj���dNBۋZ�6�F:��$����ؐ���R#;#1|����(��-���5p���9\��+�vg䛤�b,$�K���rk��V	�Dn�P
 	!+e;6_��6���ֳh�q��i*{۸C�����I|v��Ra����M��^|E����Dq8��N����7u^���q\�����~L_���0��2�k������K���E��+�ڴ��i�X���/��huӔ9�a�D$����9���� �Q���:�"vw%�<�U��>ۻʭ^-�pK;кt��?��ݗ�B�<�2��9����Ǟ�>{)VY�;�x�uMf�c�@��W�T�7�R!��Μ:��'v��6ŊߋʵZ-t���j��1t�w�V��s;�k5~$b�'�v��Ӏ��a��n��wv���RCu}x��`R����55���v"?M0��|���ޡ!��畅���;Uz�~�M���Ć�=�I�3#DO6`�۳%�"k"��7p#6#F���k�z��Ý�xǻ`�fG���҃�~�f�YE�c��W[o`rM����~Vc�4���=����J�~��	1~�V\�5	��s����PD]w��e�c
�Oǐ�1�ҧ��D�K���UO���l��;T�f>J ��p������%��,8�?H�x���e�E��ש
$
,lZ���[	���'EfW�g�ʓ�*��.S<�=B��>���:k(��^�ct�٧߰s�#��(�G.��3�-V��V�UL�.�>�8s��R�����%n��TFV/=�36���`��z���CNR% ��`A����TcC `���'aE��>�ˎ����f�9񖇊Շ���v/c⻾TYn^/7NE��@%�.Ǎm�'8��14�{�5��ٽ�yQM��cl[�Uw�E��{g���R�����t@:�q������&����:��P>T*���z�c�ݻ��t�j��2��'�&��4m�e@�3v���$-2�n�lH:Z�z;�ɨ)8Lcx��2�H��E^��(�XoȕC����]wҐ�N�)��(�����Y�d_.Dլ4)��;�|�Ԡ�v��N5�Y�%�BC�sK^,[�Y�l-__���"��
$PKg��8� Kq�Bs��!����\���� ��,vP�3[gL']�Qv< 	9��¶���,c-����1�+Až>I��J?�9��aF�R3�(��H�ּ��3��y�1|������4ZL��vN�����0/w��A;�R��E�d๴�&�R���QN��`��Y�
�{������̛e�,��4�/�!t)Y�;�,6@�F��g��N�̾;0Ֆ�(��E����D�Fވ7)ٳ`���$��$爞#,���x�aD� ����0h���ϐ=�Ur�J;�a��8׸N���u�ñ,�Z�rk������a��������ss����5����ᙱ?lf0A_����;N���'����!vx5�w�h��J)�55&}-5 ��J�'��-IN�P��9�kVL�|�]M���c�+�� �.��/r)�`��I�b�a�ʥ���n�X�h� R|����q*�1�(R��zQa�:��S��3����rt�`�ͦ"7p):Ƥ�A�ݛ�~��E�-��M<�=`���N�N�L��mR@A�Ȓ�U�}����"TZ���n6٬�rO�B�ӡ�usɣ+�e0�O
��	�As_Lb!�~j��0.����Ku�����-�9:��RA�VU}�����$V�4oJ2��l�mSS�H_1�cc~�j7�3���lG,3׺�Q^��}��ɣH=T	�!�u������;��'5��q�W�e:FN��ZS�Ol�,�n����g�ڀ2��\M�U����q�n*��B֛JQ+ʫԜ9`?6�����D�4.�9U̖��5�vn��2{� Cu��7f�,�{��5|�!f��c�Ҹ�lx>H�q�zB1�d弖�z9�:0���E���C����}(�y�'�������[�� �s����Y��:����3,Grm<�x����;tYwn�%�n
z�Q���"�u���ɭ�(��RY��1�Wx�VQ <1����?p���n�f��,G+t1��φ��|)������W���i~k�a��7�'��)h�!>o�Ƣ��'�l�-:��׾��~
�8���-�:�6�Y��a�#OC��dM�h�QM��G��3f�s�o�:�]�n��2�^��A�V(4n��vᶺ��7�5�u�ǈ�"OO����l��m�����+S? p�	�2���d�{ƘBs�]�=N�),6j�r?;.����O\�;��u=��܏`�e4��rs���AaxHy���� �X9��Og��	w��K=��� 3Z7��ڐ�l���Gh>_ӭ��8��N�P@{�\�5K�@C �S-�I^�oX�(���1��b�fN7���"��kD86J����Qd����x����e�L�ZΊ_KF7?�V��Cb��;|fV�{/�P���b�G���� �6Jg'�=��K���T��B���x�N|���Zt���ʉk�/z���TV�;�=yr�\*6����������"K�A8��<z:1J*])�jY�~����f���f��f�ܑ��&�K�{�m��e9�IU�-]�z)~JP�j���o��,&�y��G������R��;�<�k���Fk��A-t��[W�c����Z#�S��������۩�UӞ��K)��3HO���x�{�)�gY��3�n����O�]��/�%���R'����կ{ ���ԛ�@ѵ�r����2|і`��ːm�O���6>�>�h�4�]J��0�����U���,��u�� ��%0�ej�xq{U�ޠ]�9��v����`�y �x�n)�p�30s�7���?k�k�O
���{u�1-�S[jB�����}a��dz@�^�+>�ݼ�$�eG�����P:5�|N�����d�ۨ�W�g��6R���a�E��Dp)¨��C��
!�<D������k
����2��i侜��Sm%�y(q�UNլ�އ�P/+� SZ�6_����߻����2H#�p��Pg���o����Ac�P�w	as�y\2�:�� r�:K�2�&ܶiL]�=�頚w�rb4h�Փ��	������<��o"�x���Ei'�oC�Q9���$��15��?�!v2�W�	��!�^<F0O�)ɤb�G_#Ұ��6ψ, �Rֱ�N��e#{5 u�KH= ����d~S@�u( �5RB�&� �C��&�dȖ�� ݮ��O~~�9=�z�X��q���:�+�H`��WB��p �@j┲�R��I��1MĢy�6C��P^�����͟0���o�sx��1���~�ta}��MҶ�"��k���vT{5�5 �t�����16������voX���ֵJ-�^u��������@x� �)�C�&�Η��3�����'M���Q5� ?�a�QM��`�A�s��F�=$,F*�m�9�+�|���aqS�����o5iՒ����O�8~}'u�E`�I<�J;���3_���_^�W%�,K��cҜP/�sI�D!!��z�Q�F�/{j�i���.P`T�Ɓװ������Oɀ��d[����ܧ�r֞�?>£��y����׶��/|�-�����p�>7$� "�O�`�� �<c���ІԚ�]5E���)ޘ� ���> �8���_��u�@Ǔ����Ô�� �.A���n��Ζ#-�Ď��R�{��=��1��8[���z���� h��掬����*,M��3(�����⤞���&�\��{��r�Cs����j��`^˖��������x��"�ZC؀#���_��yآ��W,��mXE*ێ�w��;��r�?z��E��i�y�)�%�'���*����S��T���F����O�Y�q�E���fDqû�h� �d�2��UH�~e���{���׀��8.Z��5�L�YD��a�@�b��(�H�l�:��=0�#jאY��4�l���N1n���e�{	�n6L�}Y��{�������{0
Ţ�7�\��Gv�(�8T�X�\.�g�`��56��	�ӛ�����"x��x�W͝k1��b/>nMw���>!p�/�4|A~e�&�R�lǊ��/sʵ$�n��H�q���^�"d�R{�L�!�<����kS��.�8o�M�%6�5K�����C���[�kS�!��#��k+�2װ�ٓ�!���7Y�*0|#ڹ^6�'PlG��+9��%&�3f6m���=^tn��(Uz�X��=�ǝO��S��*���,�f1�m=�$ /��;�7����q��c��Y6���i�#��t��>�lE5V���ʵ�"�f��ʇ�����S�x�W�d^=�ӽ��`����B����iŤ�P�K�Y$S=	"����jH��-0s2V
)o�SB�G��A�K��8e�L�]� �;W��Q�}J��Cl6+"�_��n�g"OE���lx����8��Tӕs�jPr!;z�pX41����{Ql����ͪN�'��l��3�����.��:,޼�AH �ޘ%�j��N�1�] �?�3�e�3���.�� o�y�̧<D~����Ա��V��rŹ����I,��N0�v��֍����V].o�v�hr
�x����ϱ�;���Gb��y"�Zg�&o'0E�8hD~S��Hy�V�S�#J��1�-T��;�v?���:o �?3q�ǫY����N6X?�VQ�s�O;
�*�o5Dg $�xtw��O�(���h;
��*!�K��C���d��^�o��N�2��L�:����;h-CP�[���jhL�o��.8z��@��*�<%7��RvP,5Ӥ�%.6���R� F�;��(�!FW����j���4e��d�E����I�ǃ:�W8���:O�pf�<L��=�=+U�u�K`�O�������g���n2�����8&>��k΅x��(hcZ �G�6^��4�R?l�î�)�~'��AX���� �l�=x�%7�Z���2mQ�G֩eW��8#������ʃe�p�6øē��N�QӍ1f��5���F�b�V�Ht٧]nb���hL�Z{�����d��y����C�ȂRsKbR�'���o%�B��b��e!����,	�zVU4�$�k^���j��B]��'z�&����j����������L�!n��T�)H�HF�v)���&�俢U�'�|_���i�t�d���I��1;Wxܖ�Y=(L.�k��)|?0�22B��Dz����&`����:���H�	Ƒ9
� ��y���S%���3ne,�{��,ǒ`&��j.�R����Zi�?�!Sm�O
�]u�0j���$����!��XtD_ؽ�����rT?�n8����D�����{U?�(��׷M["����Ʈߡ@DU�& �(j�n����Gi�<%�>����Oߌ�ok3崂�'��a���������Yxu����7�o�Z�y,�<�C�A�8Uao�H6S�1Y�dh���a�	�Ƨ�gׁA�D�e+?i�rX�8�*�Ƴ1�w��s�&�n��8<J�mƤ���߆�5�����2�>�
��e����g�Ɔ!r�N\�mo"�zM�_��5SF�_zY���r����7�]?y��������$���+4�;"��L������H�gkƥ��(������;3Mi��M)͛�+7
����@ο���U�_����c���W��3�/�4�n?k{��5�pt����/��v�^~��@��m*˩�(�!)0!�6~r��=g����뭡}g�tP�u��H���v�����|.TGX@ؗ[��[�u�#e�i�*焑
�7ht��4%zIa֘���"�sM
3�p����I�g��mי��<O^4���9�E��&O�(x�+���R5�F}��w�+h��W΃ֻΘ��T���W��
E�4�F!��t^Y��`ٟN�h�ŝ��Rs���d��,IU2���k|~k�i���Y��}�ly2@��!��X�����f��RO,��;�7�mѺ�vTT]N2��I�s�v�Mϕ�	�~�,�K��`��Z�y�|e\]��:��� b,�P�dM�&l_�"|�uj"W�E��(9|�?gL}/�:dZ�����c�ph�x��4i_8Z�+��Pq�g��h|%�}ld|����Blo6-)���ܸT�Ï�_�:HNCi�s���ĪpB���0&\��cP��R��F�O"
E�Nd�T H�3�7��O�H�<LBꏙ�R��L�Ǉ	�i6��%���)fja��$1���� ���S\>h�|�R�RqGD�0ΙUq�U��ܒ��4�^C�%��x��﵊>�\�]���UѝA�&�})OH�x�)��no*w�#`$?4X��߰�3���Q/�z�EwE'�ed��ng~�?ړ�N�<��#S�/�w�[�z�,��m��/:���Y�8"�'	��(�����rظ-�CoEhi~���I��iGs������A���$わ�J����~���Ċٹ����r�-�q��rHŨҹ������k��9l����ڙ��FDS�4����I��X�z#؇��k�`�Oᬚ&��&x�p?�ڲ�
�G~t�4���a&,��܊p�����B؄���}�b㴨.{��y�f����@`%��9>�
�Z����*���sp�� ��`�n�G�z�&�x���q��|���\������@2K�kX� Wa�A�N@&{9a४������!ec?=�1D䪶,��]Qt��b��נ��5�0z�Sܥ�E�ԟ'�[�p��<^?(=�ҙ��bĪ��۴U�S�9V�����o4w}�F�h��w��ovu� ������mP������
�"g><|Sv�߂�U����-�ծ���s����Kϋ�6�N�~)˜?h�>=���-P�Ċ�>҃b.	�k��8�4��&�yh�!��8�t���J��;u�ȵ#d~>p7��o���{~�f�Z�ip�T�f ��w���ղj�j�>p@����y=��b*�'CU�GB�\ni�N���OIsB�K��L�hɭh�G�/*T�[6�mS���#Z��^��	>��]h�s�x�0�L�ǎ�JBl���:���'RDz�&fz;9 ܴUf��l��Q�E� 5* A%�}��? �s	T�� ~�T3?ڪ�i�ssK҄������;�}?�d���b�U� n����p�Y'�;����N�����"߸V�3UM�<�9ݝy�Jf��b�dL#�`�1������|�q@:0b~��~�9��M5���d��Jb�P�� ����ш��4�d-��(O*zV�O%m�\51;����􊳼}���n*9�T[���p�-��G�٫>,	b��Ox�O�e"�ϴ1h�6�#�
��*L����g�=��<(i�j������ D�r�oGf��q���j��V%oN��`*F ��,��D"���/�Pc�Tu�'��1��M�!��^�D�)��3"竉+�F`�l��fh��o`�e�~|�xE1Č�:r��c����[Q��;�iM2��n,� �����&�
� ��X�*��w;kG�U�=�r(�]����2����%9fN��Nf��y6w�NםȨ4�@�S�Ǽ�?f����Pwv��{�:ة"�-5�>������7�������#�w?AX9�?��x���Ь��t�p����^8�i�h�Qd�hlK��E��4�'*G9�9�o/����gpyަ�����6oDPIm#�h�I|��N�Tl@
���d���u�%5��w��S����SxX��E�W.���s w��H)�]�j���P�.S�^��J�$�*d!_�Bǫ��(�юR�k>��X��E ڹ�.�03�� �Yq���y�����瀮��F��N=��0�8K��k�(:�ˠ��%�� p����c�v�p�����)�~�vBw�w�������?^+��S���I�[�Rqzٚ�?
�=*�Met�8f���F@��/Hj!�*d�ͽ��-�wwm��?����~NB�t���ފ�wɒ,o�:�%���Ă�-f�/��Y��o��"���tv([}��:H����|��Z;��F]³##���阔�7M����:����S����U����v�H>^�ዪ�>#���*��Vȉ�� E?���]�<�!s��Q�4�@:��K�8��|���xb�dw���r�����%�'ߦ���9{9Fu�$ �ԣ�[Q��4(	?��{��ICZ�S6즂ˣs�b&��tn�O�^ ����ui���=\A3'H�)"�}aH��Q�����'1�Hf�o�.��Ӊ�����=�����������9�Oq�S+0d��=�s ��NՏ*˫�as����p6�Ӟ�?+���|��]�k�5�:-ف i0B�44q;\�0T���D�_a�;�&�\ ;W����gS����r�9�
�� '-���"a�1��6c-\��c���{q��F.��n��H������P.�Ft�s�x��.��'���I��Sk�X�5��8`����?g�h�k͔}_z�p�eBG@���̟�����`�Sp<�g<ױK��Z)�(���=9F#�u�rn�d)���1�.d��$�O?9�9)��������}G<&O��b�\P`���N��I����]�R^9"�X��Q��S�|��dh9�sf�z�$�m���~w���Db� ��Rp���s�\��I2e���?5W����a*��I�9��3�2f��a���x	��$E�r���� Go}]���S��S�=;����d�WӠ=�0�= 3ʛ��bΆ�g�^ɗS&�
���ΔN�4�����t��^�72����j�F-Ho#���C�<�iv9E���Vт�Ճ�ڔ�Q3j˓jB�!{��(�!�*,���'.����.CԎƥ�9��e��l�~-PZ����+��I��$��po9�)�l����֗8�g[�wL!�5۰�߮�r�.��^}�7x��##�đAD�����vs ��
�)�w?<a�/�o8������6R��V� 0��)�e��@Q6Q%f��
��[�?�z���������ag���e���IGu��c��˨5Pw�X�P�P��1g㙿g8I�+?���X6�llw�Gu�O�����ڴ#ްd��U{+���a��m��I�eP^�(M�6�6b�P�ܳ�+��0WeG�~X��H�<�E�b:�6J^-J:N�:� �D��a���qɞ����Ԭ��?%P���(�ۗXY�+�]�<y=A�D�S�<�m�F8j��	�ӏ��=�b�#w�(qh o�����m���<�0�@����CQ�َ7rLn�������\���ى旋�E�w�{���@�S�V.��{^����zP�8�3K�AS�	Q
K��:��8�4@î�l�W7��A�60l����^k�0t(M0_q�V�O����X�?n������@Τ�X$N��!ݰv9g[��.�#$�Z��~UۀN��$����ɛʫ���J&�5a��%eo�%��ۯ&��6L<sO�d͜<L1®���)~<�����C	kɤ"D#���MB������Әd������:��ўJ�6��I�Hi!��1�<�@�^qIi�	C#ҳZH��m�x>zh��H�>�����
*^¹�����f_�*��#�$W���r|.��M0��T��)��E�"�Fz����ƋR�	����������=�Uz���m���F��(>E����*zna�Q�X��$ޱ��w�AM�AK0�fY-�D������w��jd�!��]�� �I�`��U�#���ѭ�������+q.96蹑���7�r��ߐ1$�1c��v���Qm�_Ǳh#�3�c���`�3Oݨo�Աϭa<���	 `cxZ��- ����,�=����#�dLaӝ~�i/ӟ���[��-�I�>T�*��ej����΄!��3���X�.��Ow{S����+���F4�ʊ�u���F8n�#�ΰ=��n��%"n��@�:Ƚ�;�� ��	����?�y*�VR-�t7k�R�u�C�)��I�N��S�T��>>����p:��5'�"�
r�=Xe�:z����"s7##e��H�K�ҿ�#��fhKҺ6�Uעv"Z� "��Oߏ �4�DD�-�ҒW�۾�O�d	�1ט�g��EhX��Ie:C!�3�P�j"貨�f�I�|ܣ��3iT��ih����<�R��-�ZrP@hX�G��A�C�y+G�7�6j����� ������1eŠ�LL*��o�~�m	�p$y���ܩ��:�e.j���'��@{45���#���8{c<@k͆���f�[���B�8F����GoV�rEz�,��:������y :�ob.��F�T�C?�����\Ee��و��٢��3��"e.���X�|;W4<�P$]n�6��|*(92���h�?A�����l�-i����h����[�OZ�sq�N��qc���g�qI��>���p	�ƶf�e�Y���['�4iyudд�|b���3	���÷W0�"��FGf]��?�Ue0�[΀��Td�(F��|
}�lXDw[��_��k�U�Z�k�`f
(�ju�.�1�I��dz�qʊ�S��ICE�_d�lz�GcD��y���NϷ��$e� * S�8�Z(�L�$H���kC/��� dҷf*�J���ձ�|r����Y�@���0HQg1!��iA�K��Q��b�1��148'���T1��яmQ��1Y�,s��E�0��>�]N���F�L��9ԩWE�d�YҞ�!��}�<<��ʚ�e]�?P��C�F�i�O���)�e�����d<3���3���%�/�/A*�i{����U�-���5	d^��}����m�������R����G�_
��[J'�I��*]�����{�_�#��$�VB��t��5�gnml9-�^R��1��KtT��z�p�E�0v	j�tǣ�������I�GLa����7w��0ـ7i=�,��7���Z�=*��5��G%��_�d/޶�]�=�9�� `{2�L�X4*�����D������n'�,<8�m?m6ad&���j��X���������h���w�_�1#s�W�|���XU��j'ëT���������G��1��k,z��r2m'D@��|�?�+{��(F�|�k���D�.Zh4�{�;e��@y��x���A�F@��:��ާ����hA��.���E_/��`B���g����X�K���Le�YXM�G��2��~� X�P��ݜ+��N����᩟|�g�f^��`�������
jaswy��\����\����C��M^|ߝ�
/9�+�5����C��L4?5��[p\�ҮZX�>Qzr���҅�-޺UqO͡���?m��o��hD��~�����`�Yt<�w}a,������ZU{CJ�_&5����%��:B?ϑ�����|����c?�]�$�n���z@j=����+2�S��/�2�Ғ����'�vW������!5�m #� 6��]D6���ngG����X.��ʼ$�|�8���zȏ}�]i*=���@&��ݸ��F˄:8�hJ���mߚlIg�F���ZF`���'�>��vͷGI�܊�Ө��L��9�x9��'��A��dq%ni����q�fI0<�j�F����E�P&�S���~xA���~2Cᙵd���[`�z��K;�ً)��#D)mä�N��ܪ��4Z����ϧ*�K�3
ʸg6?�)ݬOyr�*�X�F�5�	 �D7�csvJ�ii>V$X��Wx������M3N4ǥ�ܯ���� �y3�y"�9*��0���h�����9֞�A���Fy�����Hy@{3�\��
�x8�,J8�iՏ�:e��1��5zQ��f��}�g�%�0�=Z���X�X�/fCc�)��f��$�:�+$�~ ��P�C��V �)f�LUT�bq>8$�]@]P(�_����I����MB��Y*@��szv�cb��jb�$�����~����a�T��V��x��I� cn�$ڶdB�ct�c�zM�<xU�ucݯ�M���@#jN>ʷ<��n7�a�����>�:���JV(���(�v�]ME.(�:`4����P�%�ZN67���+�oXZ�\4�[�k��/p����t��sS �I��J�Pa��6ɧNdB�|=�4���/k�A�^���	D�����N ~YqSu�p�@�\h��eh1cU��hI="��8_8�����%�e}�T��j�ܒc��4��6��픶��k/�h�7z��M1���%���`緓՚x�|WzU�զ]0Q�A{���(�Q虅Bթ���|�0�\/�.�����x��]�14͹�K	3�#��V�<_�J�ج:"�"�RV�ɸ*9V�0u��wS^:�hh��`M�%��KK�{!},�͇&6���
�˶-��a�'�ag�YS_�$���l�|��\)�gT��?��JIH��7p,��Q���:��Z#��tJ�,��ATI�Sfᆍ�ɫ]?�%8䨍I��k����J�m�^j�^S�Zd%�
���|��7����8lS���٫h�OԒ$�:M^	�'���k@����6�>wy�5�kF�Q)��b�S�Y$�O�o�&CP�>r�s�bx�t�*r��>U���d�Q~a�r|��HN���Q/�%��.��&f��YT�y����֒!5����{��zH. ��a~大3紿��A-��҅��9)m�HVO}�ɿA"�&���U���9`:wh�%b��^����Wq9F�AZ�eQg`����SK���mՎ�"��6�&};yR���[bA��2J��X2rV��fz>�u.шn�?��?pEٕF,�i蜯7��q>ʛ�! �����	����1�����wS������f͖������F�r����4y�WP�}�>��'�7#�$�:� �0�
ܗ�R��!3��;�V���n��1�?�/C4?�}|���d���W��[�6�i5�A���.���>2B��5��H� ���қ�Q��ڌ9�j�DH�J���U�l���-T�nm��ݦ+�MV�F'��:�v�@�s8�±5i�'��إW�������+��؆c��/0(�N>��ȗ�"�3l�K�T�����B�Mv.a6����3?��֨9�0�L$���\.H�V.d��u�d�/��NIt�a���V��h�طo���1"@�B��N��H�9^r;
l��<��l-V�o=���gs�g>��������d�4�_cɛOa-L2vP��5���Z��r(VV�H`�65��	��d-�����T�˥kkiLy0�&��[��كl��,�F��EPS�p�`�3��B�i
l�������?)�{��Ņ�B�t#j�!%���&���������nA�S��0�����!���Z4icQG��bk��Z�JE���C���e�s��yq�]�2>�!��l��Qbt��R���>�kNk΅�Y\sk���"��m<�%�!H��[m��|�yDBi:$hZ
$��5�"͚}�g�5��w:���D��	s���"������wjb>J���u�,��M����8"*�	����
�/L��!c*�)�nf���H�%�9�"λY����~p�����Y㩰��c<-a�H�l���T�(N��@��j"pMԖ���句(;�IG_Dh���c_.��f��!��'�^�����<�>�8HL�W�e��-�2�Vu�����Э�j
������?-j����`� �eh����N�lo�����ا2&�m��fEk{�=�� yAB\9#
�;:�w�G�<��,��kߵ��J\~&�߲S�1�\n�N[sO�ؕ���'-��:F�1���rx�ڠ�.U�]���;\ ��Nq�o%n!���"�A��O�m��_ts����FY2#Z����}�Ax��]�LQ�K�w>������d��l��4;�UC�l��F��rG5��X菘Q�p��tQh��	�F4��`0y">�9HN4��P�E5�VW�ѥ�:5oL2��]�x���{�^�fC���TI���l�����|G��DH�+��ί]�
$^j;U~~�ު��[	4u���մ+^?)v[��))0Z��l���iiVm/{Ʋ�Դ��"��>8�Yh�O��2&[l�v4�+{k<�s��&�n��gFj�"�B�y��O�\`�H^-v�`�]�]�#��:��6�2���<aS7k���+b(�TY�Ś8�W�K8���Oa6*�e�a�kF�辖��V
�hJ4�L��	W��|�;��L:�K�ʈ0��M3
�c֛�b����m�%�xQ,��>7���̚ڮ6���15�O $K�8���* ��Q*c�j���9^C�Z�o}������w�#��1C�n�X�#hl�̧�m��?����yX������vg�������Ͷ��\N_�B�Q�KN�"/U�����{=�ҟ�9-�E����m��[����������K)׫5�w�c���M5nE\�ָ�Sɿ��Ln41>��4�ǯ�AvC�
K��4Y�^W��H�[��J�)J��Z��;��o���>(!'��nI���Z�٬���E�Yqڃ����ok����j	NM��8;�7���v�P�.�.[�#h	7�E0�����V%���!k�T\�#A,VXB��������aN�z|V�B��p��#Áa��x�_�_v���bg�䩀�M-'�涢É�t�3�y�F͜Mη?�+��#pH�.K�c�l)�峨��bEo�o��ċ���.j�!�ä]،�Z�z���b�߫I� ��J码5Ăe���ϒ�FEpv���:2�nW��Ь��|*���q<����f�zQ.ٳL��~X���c���b����T�eאX}d�A���4O�zo+d?z?8��+��6��_y�s�ɰa�z&�I�H/#,Wǣ��I��9ei`"�g�Q�`1Tb�f76�'���;�H~%�qvh�F5�����jr<3�b�0{�r��e�Bt_^�����˶�T83��ӓ#r!�[����ˑ´?=�V+Y��:zr5ݲ��÷��N�T)O��H�O)A��7)�g���zTE��1�F�pQZ�u)�
��_�����Os̻�Z�-�P/gP�����$��zp�:��a��T{�Ν��:*}�GR�)̖��jv�a���c華�"�B�dF�N�7w!<���FIA�J0�����9U:�Ln�6㼺�o*���g��\u	Oh���3�ň�}�Q�#����0F�[��cX�G8
�\���u�Mk���t��qU�a9��C��':��&��>©�q��.V����|S`+`z8�\��{�,LqO�7�P����N�
ޡŰX�;��_ϻ�s�.�k'oT5�����+�!|���)�q��\�0�5�$�����Y�E�d �u�d�%V��%g�Ĉ���K�_��.C�ʅt/X��n�f.MA��0娡��X"�Z�PD��J�+s������B��xwZy\�2G}d�nje���-@z�1�l��$Hvh������V�cP�6��Y��P���f�Ӯ@�����Jon7n"r��W0P�Vg��FHNz�]b������ǻ;�!1r9:T��i���N#|F���Qg=���?0�:�$��7���Yt��kk�M*���نD��1�,��d���_W��?d�#��mq�R���O��	�t7_��A�`��5K��V`��`�SbP�W`�.оjw�ew���8�i8B��S8�
v��bl6�kf�Av?ճ8 �c(�̴\۠|��.�5��r�ɮ�|r�Su^Fuo���
�o�{2t��U�w
��=��q���,E5�*�X5�0ݦ�4C|*����C������i�$�<�笥�-���d���5�I�F�qX��4�hI@���Ǟ"�Chf�H���E������(�6��CeI����G���	j=?a��&����u��sa�w�o�)��nˍ�܈'�t�f),ZR{��M�Ȧ��$�����/������,RRgI�Z��-� ����4&����NF����uy-��z	��k�� G�\�hTc��/4�^�&��g"pYV}fa;��Ù%�wk~Ꝑ-UC8B��Լ7Diw��n�3�V������c��ڌ�v��ށ�'5�;Ǆ����ok��􄁹�t�3�q�~�T�]`�>t�p�tv�D�R�b�J�M��w�6�)4Z%!Kok�T��_�s��қ����`14{_��Z����rT��f��`�&���<�XW�/@������.�~���b7f<̚��C5��P�4����u�Ң�r]�V��Ǐ$0��pt{,���q}��xIMj�X��o\B|N�؄��]tΠ*���o��z�.��i��u�噮3S;�ѿ�ӌw*���쌷v�m��fkb����1���M	�F�A�t�K���7���2 �?<iKg:�O�[�,�]�"��T=�ҶL(�}1O{�HލV@��+9�l�U�KpYf�E¯iu���9i��=L�.�G��0<KdWG�(R��ڌ>��ha7Z��sz�)���NA���]�*]/��f�W�����&c\�����C�
f� �$9b�%|и1a�����˞�v	�6�P5j��*=r~dV�(x�[����//qd�_Iq�^W�J�<�~���d�b�'�:C��Ȉ��S��)Y޺<�?f2���;O����r�k���"��u� N��XZA�c�@Dl�o���U�9o����9�SY��+M|@��Pv��-�j�#�D}p4�&ے���?�es�9��{����w<a�ƾ�#�)���E	��N�Y�}���d��e��x�qW�ؓ��ES3�-��K !Shj|H�W����υ���T��VD��8�m1�->�M�5��\��yA/�'c���n��Y"T���œ6B�= y]�q�ڸ�"h���^T�YF1�s��dHa�e�2��6m'$�;7��<X�M�fZ_���O�>�B��\7��V ]}�i�ӭ��
�Z?�C�ER���9<&�o�1���W��A��g��c_t�DXC�e���W�|����3��%~�v^�/��LBwg�ի�5W�7-?��E��@/z��ؕ�d�����mЌ��@-��&h��FTv�Q��I���89�L�_����0M�8�0����$o��=��0 �V���=����z	x'�G��<�����v�b��{T�E�Sx�J�!G�j�[�,�WׂrYf�����ǈx�g�6~E.Jxܯ��_����!2�\&�*�2������-��;-�*�x�A_�2��<�L�	��B���f���}՘��6����v_��FjB�8]����^RX�>Z��-ߦ����_+�B%�X�I�i��fD�<�g�6��?�὎��*[^V?��C!~��r*�j���4u?���^�b����Hj�c31����Α�N+�r����.Z�����;��껑.�!$���޺8wP�uUsk�Cφk�m�*+��c�����
�@�7��f*1bQƫqy��Q�п�I���~�Hjd��(����|cd���	K�X�H៹	+j����Fh��ޤ�����R�������)�X]a ��ac�n\�{��`����0���7�֋qI���qE�<6�����̲�����᫟�=����x���v3��^o�9�޻4�C�>��*W�f��^ۙ�wQ���_;R���o��rG�J	�;WX��(o� zt���D�&�x�
!��!��]n��o����mq��X��,��Ѭ��A�j�W����/��.��ܵ�T��.s�4�
�ڊF���_�M`�S���ƅ���}�t�����=9��5+X�s�%����Vmp�䰦�	����!�oΨ�9	Sfq��I䎥�lA|�O��i�B���E��Yoc��m����#"L2�$�l���
~��a'T~�jG�5��N�:;m}c+�ag���b��C�2y�Û/Y-�ӯ�Y�2(�Ӌ5�5h����-'^ߒ���GxOR5&�t#��ss�=D���1�N�X_2>���H2��\T+mWB�oF��B^n�2_e������}�=�B4R�sq!t[W��;� ��|F
�=���r89fX��Or��I�����B xrZ�?z >�6��<n.�]9ᶀP�D�+�^��{׃M9�!Ě�������g�+�u��*�-�^�_���(9�O������h�<WG�] ���~T�j�'���v��Ku���k���oVgUL.>ӫO��I��s_;��]yyv(��]�F�~�)�����A�e�H�x�J��q�̫��� n�2�#��;�����{���¡��!��������݅��,�s���)����Oa8X�v���ʿ[�����<>ۑ�}�v�`>�w�� ��ާ��/e�F	ݷ�ϴ��\GP}�dW5��9B�w�?I����	��'h9d�Gi1����a���-`����)<5_97m�س���n�di����Н?ߧ�o�g���_d�����32.�R�2@�=t����U5gE����V����|��f0��K������p��e>�-���"h�C��p8ĥ/��lJ@ȟ����I#�"�߾�/�t��}3p��A썮&��c���Zr�7Yo ��4�H���J�.:&�u2�9�4��{萤�=o��t�mr��i�`�!Wb�����Z�/��#���wȇ|\ĨQ���]?;	<����Ոx�r��"3�:�o������>R:���5
��U��+ir�h���|�?��ۭ=$~O%RE�VJw��Ms�r3�k��}�-����]��1�
n�`�x�����+k�jA!$�9h����V$.LYUU����,<jfn�V����)9R(b�1��8�g8+��/�-��¡���/���/�����G&�����+����g�%�������a�Ұ�O��
^�'�e^&��*���Uq_D��X7?G�=�Ty�O��}�,|R�TQ?�(��V�g:	rՅL�=���=I��\�-�
K�������[Y�=���kS�L՛�Tc�7�g��L;<#=и} ������~��.i����4f���s�Z�'��ǗIK\%�!@p�AШ�iAj5���2,�ӝ��]#2�^�fy����:��fڵ�d�'8���m��DS�S�{��Gآ !k�����P$S�D}j7��m���e�艔u���2.2����X���!x+Dz-���G�L��W��߆��h�|e��;ci�X�����dS�Ův�x�j5�H�R>���6��I �vpZ� �f3�2h�^�ܠ��NNTN�^���w����v'd�}I��4Blt���6�	���gN�4_F���_�����C�"V*�#������n�/��=aLP3c�e���k�M���x��g��4��K-#y�(m�,f��ƏY8�o��x!�E��1�:K�L��	)%���EMM�^fC\r��������y���c�`n��r���r��)5���R`Ck|A�4�y	�Q�# u�/�4�B:X��?� ;(� t�Y���\��PlŁ��ǃ$S��{�����K�g'U�u_�4)�c�ccQ޴@�]�w
���&�J�tuHQ'KZw��%���^4����*��Y��:�v@�i���ʩm�ޘ�<���
�^+���N �mpD��W��\��n��jb��(\�
���j��.��vP{ ���g���>�l�1�~��ӆ F�[�lɭ-�*��F��Ǚ�\�.Jꕣ	P�UE��\6�v`�?;��FX�5UM��\I^�'��V�¶G*�2���wΈ�0y��+�<O����ƴ5��\uo��FYz��Oq%�tUz�ml���a��� R1������׫A�3� ^�2��(/B�!�N ��!�X���g0=��D�g��?��������/{7a
�K�K��m�;/Ű1VB���������QD��<E�Z�$�[6<'�KP�����;��n��56��}u����&>4#�ɺY�+����v8nW���V��g����_�<��/�^v�>��I�}�=����� ?��G�������粞��nʃa"�1x<�K4g��V�lH�@�*
d�5a����5�kT���,�%,��6�M�< :)Ԥk��?�n�`������s_���,�"��߆�&0?�ȹ� �����Z������q�EIN@��O�(2�R�;I�#i7��%�����Sl��^�B�/��J��+���'����R~�o��Q�6`�� 2��`׃%.Y����_jj<h��.T��\���ֽ��/)��e-����n6ɒ�5<����l����Y�60v���G{���B�����!�wg��>EHvS����]&���n�	��)��|�e��H���ߘ���A?_B����H\����I3��"�}�����hrc�������"�f�f@\������!y���4�4�	x�CNX[4�6��m�5DX�p�ʔ�0���]�×(�ԹV�y�Z��f��E`��5�&�.�dtg�Fq�����'��fox9o�J��\NZ�q+���W���4a2�h3(�h�#��؃�b��T�y��Hfv����54,�Q���<�m�#��ٱ��� ��f����k<BJ b%�S���e��V�X�#8��R��i�o:�(5{
��wX��B��9������)x_Ќ2�/za���9�-P6���Щ*��_��>.�k%Y��X�
k���԰�ל'	ѺO��M�7kg!����;��+9�?nlД�tAǆ� �ChF}СY�l"���T@�#�笄T�>K<�%�ߝ���I\<x~��8���6�ᅙ�U
�+]�72����?*�V�����c��jT�_�����M��09���˾�;����L6e�n�_yO�P���T�{J	�M���]�U�߻����Sٴ��ײ\v��E��Zf�ޟM�?D��Yx�}�CG��"CWNk�'��G(��*�#֭}�
dEEbփ��glC�|P�aKN�� �+;� �p�!�m�J���bbnܣ|"Y)	��x�]Ú[���6i|���&\�����P���Ƈ��{Mޟ��hہl.(QLR��\7��^�}g�y
���@���7�o��p-���M��ܺ^`�|I�,1�"ߴ+/�!)
��1��V_��:y�O+�'gm�`�CX�nD(+3	U���(�x¾����D�-������f-F�A�Tޚ��%����3Sq�6zd��
���h�����[��i@���I���o�s�3���珦Gc���� ���5��)�&���7�k��8ʰ$d[1�0SH��(���
L��=��0|Cv�$�눐d��&�dY6��Y�L��}6�*�[! ����M�~:��X��,t�h�\�X�(lt\<��1^-�e��������%���\D�1uG-�B�ߨ��uϳ�H��˪fW�@�➽��Tq@���������3r�I�p�[��� ~r>��KE���j�Kl�jt�B�{F%�R��x��zh����Է�j�U;���$��Ux��n4T�G .�
���O��B��\�r*����xI�͛*� {���7�B��+ӪN$��e�e��9r��6�j�����u}h1�`���n`9�-FF/���.��;e����f3�cmeK��&��T	���L<Łjw�������04�o��AU��*"���hx��`W��B�Rٔ���L�+yC�XQ�XW@���������v?�h0W6�]�-��r^�uPğ�|��y3$��v'"�B���I�0}�H��4d*�>q쥨h��$��t�ͩR�y��������s�
^��7�|�*�A�qBzB��� `l,o9������Չ��f�;K<P	9)K��4|�������<Ւ������j�	�Jت l.�t��h]?��`������r��䢰��|:H�Q�9�SY� |�^i{��?�F�@�����˿�KW���7�)b*'�����T��FD���x��?}5$����x�H��R���Kr����s��Xy����q�G�?q]��|bЌO'�R*p� �:�O�C��T���t��:��p#ߩYg{�Ty���~�M�Tʖ��*��'I�'�����T�r��C���~s��^l ұ'Ŀ�H�nM�"zEa�~�nq0z�� �4�ON�Չ���1c��r��v�%*���c���"�Ul���3���_������j��\�&�q��T"Fݺ]ܶ1fy�c�d���N����c�s�B3���)���7J��r�ԁ쪞��x�N��N���NQ�ƨ���/xت�x�蕇t�l��C��F���	[�=���V��j	�_��K!�oe'�oM���������X�a�Nρ\�y��=�Xظ�EJ��`z��tJsJ��'�'�Ty�=g�-v�ȫ�I9I����=u�DxO�7z�T8&K�z6`�6���+�1�k�qv!C^J�XŔ�P(
�-���k��1�6���XgBC�8����Y�jlkH֍��H#�e�yK�B������*�!�Nɺ�����l�w��̡�A^ˢ���!TV�D}f��Ihh/ʿ�{���k��!e���L��jzz��;HaTߨ�=�����Z���ν��+��9�4��,%�>>Y˨8 Z��u�8@ӄ�dJ���m����D~o�he���b�Мְ�mG[��-���Uv��>�±���*�u�4bI<BΤ�̻Sq�5	��=e��s�~v~�,R�̻�#9;�}Խ��S��h��PE����+O���� e%�]�����u��
�[��{�a�!P-����t��c�P��5��etCo��Cs��l�M�bJ1���*�y�w&�+��*��NU���cp^`jPv;��^8	�,9�K�)�M�������h����?&�ry��R$���J#"��ԣMYH���	�"x�{7-`�B�55��[P�@#����rF/0,]{Į������X� ��kE��|r1@Y�&	�l.Ӄ�8}�VH( ���#���,����2�>�����mx�4��V��� [La���UG�x����t��{��t����8��WB�y�V�!��+�c�#�$�eW�3\�'3�⏹&�j��*���5R�b�!=4�w�qGr����f9!�����:A��x�8�.���Q�h�;Vt�پ��^5���.k�.d�6:țX��6�o�F��E���LR��x7b�+�	��ǖK�x�;�x�#��鼗 ��5��&A�6�~�U��8������>�ߜR�G�6dP	��lǸw\h�	��E�w�bz�?��q�����;�!��-��ޫ�|���o6��{�0�f�&��20�w��@���1�_��������
�j�SSL'į�G^���ni�K D 0OnL���=�I��Ћ���8���w���G��'q�v��w�{�/�b"��Y�<��`-�+s��r�5�(A�Xޚ̂�L���Nꫥ���.)�wi����@�*����ȧ6�t7n���
[9>�`3�����tZz�S��_�pOܘ��;ہ`T1jK�e�������q�V4�2�\�x��5�Jٟ��hA�eG&��z[[�aCvI����I�R�&C2t�"׶�Ϳ;�\G�`�0�J�oyC�T�،f��E����	���Փڽ+���qN/42����Z�Z���s�
�B��0���*��m��>���-��v.��ǡ/'���`ޮQ�mI��)K�M`(M�2��{���}��.0�x�����|wX�Ҷ��f����:�Һ�Ax�? ?̢M^��<X��.WC[߃-���5)��E��ݨ�֓LW�HxT���윇[l!yoӸ���P^�'i00��?�j](v��������Ư��'���ܒu�m�P�Z�h�щ���Ĩ�}�Ai��;�>�a���H؜o��h�!<y�ĺ �
ߟ�_>�="t?�Y�~�P�`�i��5�ö�Y?���ڠ8N��R����P�i��D�_�<�:.��ɉ�+���B��,5������KGTݬ|�b�6d}Y4*E�L���W�� �8�.F�� #�G��������.c��&�T՟�`�����g���Î�_��A�ʰ��tO7�T*�D�S5�0[,�v��������ז�L��|�~��na�u/%�"�� t�(�[|�Շ����u#m���^!<�lc�X�O��Z��E�C�F�(�	y����`!-���|����i����V�ߑ_��+��ŭ��q%')lm�ɏ
!h��!~@ى�>i_ՠM�0�f&���L7�z�~�m�׽�o��08�B�ݸ�D���J�K����~�i�ĕ�v��>���Yl�2�a�𤊾���5(#٦���-Ǭ�}+���y�[�)�Z�}lW\�y���J��W�f��y��LL?�u���Y�:VF2����J��`�/�o��h�X���덻1�	n<.d��@�m(�Ɩ�t+>]��7�`2f���D*��A��*��PBX*h�ރvU�sx!�c�t�/^�E�aD9�H�ʝ�c�$��؍�#=�V�㏙���Xg���ekc�����<�(��q��t������w��6�n�H�����^�tԕf�R6��{:�����=+���x$�"� >H�V�N'$q��}�t����F0���OE8	V��!�áz�4�h=��,Zf83$�1���%����}��1�?�x�M����m��f��Jz�B����=+���;�#щ�-_��43���'��fܙ#j4��F�����YјO�K����䱫<A�v(]3�n�z��aQ���)�	ܤ��N��@_/��GC<��nO/G%�P,`�54ɐ�2A;�n�쥧��f�x��0�A�)bw�T̃����K{�5���GU��5���3r
<(~��)���Ȝs���~�չ
ʷ$��n�U�x�Y��9�>Y�R����iC1!�י��Wz���T6Ⱥf'[�/H?;4��������/�x��q���6'����e(����j���fű��L���NȊ��<8Bs��
jf�G�)���&:͹e�Y'��e;L'70F_��p!��ދ��Y��<�U��;��+Hj*���$O�D���鯌G��Ͷ7h�Y�!��h��&x�+����D��H���M��g�>�/��p�M4	���Mb�T(�8}�L��}�ߺ�D]����c���i��,�;~U~\o�4��$%ƂQ1�[߷��D�U�&�F���2�iz��.T˷����J'6�X�;-��ޅ@C(~�˰���Jɜ��v(>$�ʣ~Ϗ�h�o�Z&���	�����?�uҡn��
[`>r-S�#����:� ���u ��⮀�8��Q�!�n-��-8������J��� loX��:�]�?Q�aʇ�N�ɥ{^f��E^򺹦i����^��9}���0�����r�P��q����w
rc�`�@�WZfTd��Ǧ�&�e�!�}"}Q`v���-��O�e�O�A:��$�c���v�.Կ��E_�~�ʗ�k3u �D��-~���(ꍐ������J��aŵ̋xm�!�@�*p�ǲ��^��3`S�`��G3��O����n��zG$.a�&�a�N�����Z�]A��u�4,��b���Q���|֦+��e����@�t�9�n��{P���U��.8��r�xI�	�2�b3E�%q ��+�-�G.x�=��܊"C��q�E9��,�I���d��s���� tv�;�_����h��1��	�E����<GMcxuYH;)�X�c��iz��W[��G=e��G�q���	L"�6�:�ć#U�x�^2Ύ���B��M�'��g� �M=��f�D�=����LK��{�Bh���Bܠ���@�4��sNg�-N�����P_��%�����4��Oˊ%C ��}�+eL:Չ�A�VZ�a�S�J�pN�Q�E����~��1`�~bQ;����e���J��:T4X\�����)>�+\�底� �ȇ%���}��W�-S�^˨`'<��{����	�'�R�������p�A��CA˃��R�������j`D9%=i�'�}��z-�a?��<��;������ѕ�~�A���h�G���l���1/�ܻS2^�ZZ�U�V�ڇ��A�N��4Fx��C1�*�F��%S����M�ܼ����9�oGB���W��,�Y�� �p=�U���$�Jk��HS.�������rmc�-�-h���VW�e��·չjp,�B>�`X�<)e�>�,����Q�ƺ���m^%F�/גh�v��k�eAT�-�U.J�o����W9m�W�2�Ʈ��sguq��a{���VY'dph&�+�jp�a��7|�^��%ԛ[=o��`O����{�u�E��v����(_�]�]���Ǻq��Ҡ'�e�\��D�n��F��P��k�����&
mc·%o@Oߏ���bݖA(\��ґ#a��/�bv�]Z|����.D�Y�=Έ݌�R��Hb���1�I���a�i鯔����Ʊ'~��z����C�Q��0��R�I��dn���wu����f�ҋ��Se����ca"���ƕ���J���b������G�Sw��O����%��O��y��g�z7�h*v���B`��g�i���(<V��+��:�\��n�2=���U2���E`������< H��aA��3U��n�%�J�@����Էx��4�,368�QU�Ol��?S��b��E���#e2㚝N��Ȫ ����7@�Q��^QP<��!�5�ts�'l��w`��#~���!ԟ.�Dn6���'ӤO��G0B9�%ku⫄�{�,5ɻ�=�O-�zcޑd��ey�֤o����|���up��7�f��!f��3�z��nyR��;)峑؃c�5�$�y��(���kH�l�
#���N�:>@���&ⲳz��Z��� s��߆B��_�y7|'����%f���m�%ex��z�����tl~s@]�_I��"Ĉ��iKn����;���)� "g֣Tcd�
�Ф+�R�k��[�u
��ҧ�9�u�jk����luȆ���%1���C�e�ٛn�%"n<��
{��������� �t2�}ŊN8�ۈ����ѵ�WĮ9��pc���N�dl��^�������F���ؾП�b�#���wP�*��n���9_De���}�X���@H;�����'�7�����m���m�֎m��͔�(c|67��4UE>�ZbY�O�`;
�VY*e
�x�rj5^�;���T����W	Q-F��"�������va�&9��aUSB�#��;�B����T� �]QN����ƃ�܏Y3�_O��Pi;��e��"�y��P�Wrn�c@� �c����ȴ��8
�) �?SF��+����)����d�&��M��]L����#�y1���IA�4� �ʡ3F���<�g;(r�J���j�6�SH������ڒQ�O�����mB:�o4��s�L?a�R�Cu7c���6���_!ڏçu"��<�� �|��OLD�5_���-�XJl���<bLU�g��#x�t �FF���B7���������nZ��Чn���l!w��lE��v�#�D�&���qݯ�ЅOIU	]�ʸn��.#����%�7�?��I�T�B��oS}`|3٠�����&�B-R>��������_F/���ו>�J"׬�,�5Ej#�1o4+}O��Qj��@�-ܪ�8݆��3����������i)<��I��8�zx��א0���\�9�|ߕ���Z_��e"���	
��uQB�$c~�P�O:V$���=�}`_�%�/[G�G�	�~k�w��ޜʥ:��1�z����0A��yǟ�׃����� ����1�� R�&��9ċ:A�t���^N	�e��˱H�\���De�&1�a�]-K`�G���˸��ػ��5�8��2�
Q�1����%��^��C�~���N>�`@��T��̞@�Y��ytl�˕!�wY�1�'����*=V�;���qx>B�x��3�Ԛ�L���D�Mj�'A[��e��/2��6�_��)/�D-^��m�}�lE�T(�V4��%�,�I4��9���b|�M猛f(��}g��������E*A�����01A���T���˦zɹ>�%+�����YJ�9���3"�xPܞfmL�pL5R��9�vlnѫJ�7�v_u�5>H�ŵg_�{C�[~��,Y7���{��&�o���Yif����9�'���C�L���{��Ϡ-�9����-��D��@E/��~�0�ۙ��Wc9�*~ĺ2�y��f��r:���ӧU2� 6�چ&��G*�x|ZH@��EY(�ۉc�qg�Jy�c9(H�����.��n�w���8&0��g}ަ$�/�w�o.j`'����l9?S��3ɤY��c]�.
 .4L��&�*��yn����;'�_Ѝ�� ~-J�3Ь�H}~�� ����Vm��/��C���t��3Y��oc'(���/"�r�!��)˝����A�|�#���l 5��1w��a�t��D�"p��h)����=�2�Ph�J�e�I��w̺OgV3m;��cLW�|��$�t>�m<���$nh�����g��u� �t�¸��2"4}!�9�}��K6����M�H$�\l9	f��:h���~�1�t�Da@T���7O%�O��E�E;ʽ��1�~Zj+���+�)6�D��Rᛋ��M���!�d�zX��|�e�V^�l7�2�
E9|�jYn�,����q�d�yv�CX8(�>.�H�iiZ1zDP+�L'�kg=��)�������PF?�o H��h�e�06vw�K�r0�h��ǹ%�'�u�tE�mb����I5$�z���<�N>�h���u���,��V�D7��ӥ�F�=�KZ����d2�$��)f1��Ї����	_H�Z_�ԯ�p,2ݷhu��Z4�yG��S��)U���9�-PLK�������y�l��l�l��4-�B��n����N�OA��������-�o����= !V3��޻�j�)q�
�r���[B�rz_����d}�+W�J�k(��N��v%b"�4�7.FH��kxu ���y
��x�Uhe3y�^�sً��͓h������'�2�qu�g��ꈽ"W��`S(�|�A�e���;�]bD�D���	� ��jZ��n=�v���C�z᪳D�#��ڒ�;����X�i�0���mA�P�WG)W�b4������S�J�W5��,&��w�M��+�IUV���:�Zd�V�*Y�Ο&�yycHOQ�[x�À�Ɩ�-=��I�l�KJ������J7�i�d'��:jsCk�}<���Q���TC���p�k��r�9'�'�<�<�b{��� �fQ5�'6b�`�a�n2��-9R����}�)$^T�]v�r\�nC_�P3C{��Z�g�~BBLQ�mK��RP�2�E�T���B(�k�:#0��.�'�}���c\���a� 6�o�"��1�S�q/�2[�*8&���&���Z�F�h u{��τ	`�����Y�̃������j�%�ꝸ���!PB�A�1:�؍'�ς0l��$�M���8�a�?��8 ,(飸���
IF�!�;r>@(�]��+�/���݊q�.c�?"�u�1�f��@�ax������� a�D�,B��|��B�=�k#���6��.��o�Hn2V��m�����.ߧw� �rb���t�<�[Y�$��W:����450�*�w״Kf5o9w�z'��b����B�����~C]��`�\�-g�E��!�����������'!�!�� 
�3閯Ew�W�۶�0,bC*ѧ�>�������y�FS{��A)P� ��2.�{<�0:ݬ�%�ex!��
�i��&���b*o�6��|sӨtZ����8�U[�g�J��r1�E���cAiT��t�k�K`�Uke�q������q�ì��=GXa�E�))�f�*9� !^�W3���G'��V�6���t��1�Ɇ��2�z�<�5����An��BhQ�U��R��`��W�7�h�\��A U��g6�T�/w�����g�pz�	w#��c1�_�f2�N��Zk 4 '��qZc��t
݀�RD+�">�DH���*�cMWM��_ɻԽ����3v>�{��C_��E@g��.-��ᄃ*t�lL��i�K�Ɉ���MU+�� |�6��+��
wN\D7�	�u�Xl7KD"׊���S��He�5��v7��ny8��ahBG_m�=R	����dV�d� �̈&
��<��&$;�0r�Y�J{'7�%9�@�̰W�S���ܶ��6D��u<P�2�Q�2��p1E���Ub�`��2���rv��HK�j�8�r��ґ�4�)��J�A]\��R�Ui���ݪ�}0Cc37�^��S�D寐��eŹ���J��(�*�2z��I�W�t�GJ����[����� ?���d�Ӡ��w�h�.3<����v�a�n �����6|�s�af!�Rh^6��4�lL�^����C��L#����|��叅��n���S��[w�[�s1�{�O�or�T��Dй�Ӝ����߾��m��͢��Q0z�fA%u�0s�C�a,�{Ɛ$�O�$��'c��D��~|��&����#��� �h|.��aC��l���U`��D�Y\P�N��R������g�%sd4����oU~ǵ��z��0:uE���8B�����&�1�DYE.�����z��-7�����
59�[���m���1�0Fy�����K(.;��n����:m��`����	;l@�jf"idbo��q����t�(Jx��PH��9eC�C��!�8�@R�W�h��^k?��M�0"ob������T���g�,I7Ǌxjl,�6����G��"W�Sw�>Q�7���.8����l�U<�j/U���-�Vj��w������ M �m,9��c5��@�����B�囹dy,	�o7�񕡻d+���E�Zh���N�q�	x�hO�u�)W`�7糤[��[7�T�EȈ9�a��ɼ(�Ө�#�g��v���sq�0v#Br�z��|�:���L(�v�*��H)�C^=�i��. a��]���V��ק�ۇ`�Q��պ�?�*M�hݜ?��aLOp��i�&s���2�w�+�BS�3�؊^;����.����顔��,���%��^@�������贾~ d�}���!�/v-�d���P>3���#Si8y��XNn �珋�דYPv�z̹���J@�ғ��Q�V�VmvO{����0��I)��o��m��V8e3�FT�Q�v�!�S�'V,Q5�R6�۵೤t�I��&(y,-[b��qi�ta��k�����^>�a?䏶�HT��"`���|�x*�C�������(b4�MC��;25�0�������S��k��߮l?���˜�}��c���7��}�{��N �#}�I����lq$�^���y��n�:�T� �LD�rڇ	'i~�IPkVwa���+�;A���s����V��F��R<�;]"��]��"�r@<5MMJ�ϖ�˞�2�f����-F'�}O[`j<uhE��P<xl{b��{�&&y�o��ݧ-,�d:Ϭ&���z�smj��$7р����� 7�ׁR@���F���-¤  QH`�'U1�H-� V¢������t+���`"��f�5�"�z$�耧�=���[���ǩ7��&P����:�|R��v�hRt�JD��b?UǄ]�1���M��ܓ��d�}op�ȕ��?#�Ԏ����Ɩ���P2 ������_����1D��!���w����u��$��	��K��3���h
xc#L@>�/_���>��?)2�FQ�r��'R��tH���x�H8΂��Q��i4�4�Z^3z�G�R�:NB���8d�t7/�#�`��#Α|P��<�z��!`�zWY�!�|z�����q6PT�T�ӕ��Ͳ�e�ɗz�0rv1�O�P@�,lv�,,+����������͎�i�@�tk���:3,R���ά��'x�?��Ǧ��M�������ͻ��A��+&en�
-��',�9�w�'f�܉��4�T��Rs�I���뵚rY,.�����t��F#��72y�Q��A�[")_� "7ɂ���f��G O�>B�T߽e����˱�K��������aRn����RF��1&2!�|rcƬ��K�Uh�L�9+�>r�9q����
.���V9���E�����������Vl�ka�<z,�3�0�\���K�i;�P��:蚥.Ae*Rf*������bF�ݷ�"��U���^~�<�2�;�KWe�;z{|����Eqm��:%��X��Q��������K����J�3**c���� /��J�`�����kqF�7T2�#XZOǁ��~(ۮ�^qL��їm�|��o���W��hi�P}T席�Txl�g��LȞczG�1���?����tkG��"C42<�I�D9)_c������K�x�pj
t_�96m��o�,�1��&��;�g�
����w�]�l�?1&���� +�T;-Y�+�TԀ;�G/΂`�����~l�2Aٌ�Sf�Q���P����s�1B�1�_�F�P�[ �������#ŠG��?NU�*���F3r�8J�:A+�F��	yt�޵o:�<��88φ)nz�Q!��.�-��y@�ގR.-x�6�y����>��'m��̓#ЉĨ ��<ko]K	[j��D��Aʧ��=�y�s;�hQX]1� ��a��ᙨPfYĊ;@Q)��boc'��<ٸ!uyW(�$�4.H�������AO[�}�&Lh�0�6�62���	$���T��D�H�X�;�n�}OEt"֭���FR{��F]��æ��R*b(��m`�)SnTp)L^����.�I��������sb[�3&I��]����Zw�y�h�e��X0����ۯb���X���ݕ_6��c>�	� y�_�ћ�;RY���D�f� <M{�	�~�hu�������l�)Ҵg.�xNi���#O���Ԡ�zh��|��䯖uG.~C]��FG�8t)N&��v���4:J|�����+y������$8��*�?�qC�g����*�M�[�(�Z�S�N���蛼#]Zp��H5���y���8����#����R�,oQ���o�6#�y�+lݹ�҄~OnY��Ƭ^5SK��C��cK
ҐDf&8�)	b̺p+c�i�q?���
E�yN�@'KΚ0>�;^�em [�.b�}&8�ۂ1Oj�3ؠ�&��T>���G��LH�y�ڼ���(�����xV=��7b��J�u�c�2K��`}�<�,���_����� ]�,�.7S^$���DH3�@��zN��|�i��6��З!�E �z��H1�{h7�w=�h\�	�C�
%� ��<����z'r*�'3�0�~�'����>�^�]3
T�?&�°jRhm�t�{��x�f8�j�r�Xz��Td���;}Ld��.���$���8N�R����E�Ѝ�����l��Oi�����u��{��R:��3�rL����>8G�N4ɸ������ږ~��´����P�|8�""�	�^Uo5����=QR8n�T��'o@��%o+��7��G�T�l;�}�#��kT���K?�\�=Mq��p`�h���A�L�]�
3:^��Z�$P� ��v��j �ڴ2���$@���}�0 �_n�W���ve݊���b�X5;2]�r.�I����Z�(@���(���ڍ:����O(g6�d6��=%=�3�ou�7ޏC��P�����������D+ y1u��j$j��n?��0W���t�Bʅ�I��Kxn&�oթ ��#��򢮉D6�%� =�ZŦ'f�ֹ�?���˦����P�l�\���n�9����ۊiWR9�����ɭ$�v�C'T��6��6�'�b%�Z}�XO�E��j��P��������q�(�R��Nє=H�l=�f+���̩���{hQr��9D�?k���0��WeM��&�G�ƙ��re���z$��"��V9���թ�D�#����̂i��k�B25��½�L��T��l�������A�)�LP�����"�e^
�f�G��˅#]�Lg��D�N]�j�ڦs��E�P�54�-�w�K��VD���Q��
�7ࠏ�w�Z��O /cn��[Ԙ�1Usrg���1��^�Z�����굇Qĵ���Q"��=}���^|����h��V�~��������=�*f,�A�K(�95+��wm�:�� �N�QZ�А�݊�Y�+xI�HBJ4������&G�Q(����?y�D�ʠ�I�1���_OV�x"Mw��k�"mh��F��Z +�6El��>Mu�=%�G�\z�Wݸb����GL�x���5{���Dnd��e(��:dT���8�E#G�Y�I/|_�o��MO������������8�e|����ePӾE�_Vz��>��E����-O%��ѐ�˥�P�G���[�U�=�!��O�Bj���*��J��s�� [���e� >jf%#B�n��Bzb��7�{��&O97Ƶ����;.pgy>������*<�O?I��i6�ί�ðF��+�'�p�;�Ddɟ�z�8�~	������i�R�����*�Rp]�N����(��I�x�����~�E��Th�Ǌ�δ��R~m�s�׏s��&D]a�][	�>=�B!�}���P�I�$[�A#�Vy=U���]������:Be��1�[Pi#6.#L�fR�0x����\����H�GR��U⋢����8��W�e,BLyy7�>+�v���w�`�t��:���p'՛'"�;5��&���۟�p5���4� �@Y�?�ONUMl�q�6����7؈�*n�CQ��8V�L�9�Tc,�Ί���ޛ>�	Ö��[�J��n�hŽ���3{Ys���]����(��s�4~%�������Uj��GM)�>�����e��^�J��AJ^o�Fܣ�U㞺���)hΉK�:;��y�'m3���SE�t�#��)�o�j�@�3F��x,�ӕ��;�Bv�y��	��1��5�,�uXY�)�(�ĉ'���[�%=�8������+(�f?����u��^`e3#Y^��*k�A�^���FF^[�q[s}�uo�w����Cn�1���*� �.5�:#z�|]���"��I���'�f�����~3@�<��ʖ�V+M��n_����~,1��>�z��Oy!j!��Ҭ��p�Ka���u��+SH�BQ#�I�rd�����YI�',�*�tF�ᦞ�(/\?��%!���t�(3g����jݛ�Q/	U�VxYUư�3&t�X��#f�K��4�^T�j�p;-�IO�4�<Q��Q����b����R�Q9;�J�>+y�Pu�����D���1cB�Y��0�@`t��|����J�)��\�:<RChX����yt��;L(��=Fc�0�lŻ�֣��:��)�ڹ�9�Q˲+��	�T����zXF��53�x@���A&��酨�%�4�ƽj>�͑� ��x�����t��O��o�Dԛ4����c�@����O���*;��o�mN��VO�kc5��>9݇o<*�9��p��.k"R2���&d8r�x(��tޟ�3ST?��F��e�8���]Ʀ�,��'_�4EM�n'T��%��?j<��㵬Cà���EaoW���b��4HX�rz-�}�WU�HFK�|p)~Z�� ��u�|�fb��2Ԩ�1��7�e����J���-����k =�؟dK�"��$����uVR�J�G�_m��	�M���󰁃�ig�[g�=M��1e��9�:�Na�;gԆ���M��t���B���`���`m�M�̯�T7~]�ͱ��U@�D ��++��|�-�-�(ց�9p�~�eQC��эݥ"�݅O���]Ch?���Ğ��*�~��&2��jwX��ZR=RX��W���)��C��\�K��g@�@-2��b�[#����(A���1���
W:Y�}��L������/�D[���,9B-L��܏-ad�܇vR�Z��*�Ek|�\�;�ڍx�49Y(�Y�9B�"(+�*#~0l�܀QB�� ڏ����D���#N5
�|!�>�d�:�=_ٽs	�&���E�8Y�D�0~n�'jIS
ugY���g�\�2<��$ӯ9�ĵ(Ύ������-�5��׀!�c��R��Q�����47O8����W���q+�"T�,/a'}�7glYDn&�������l߸{����+A���gs�R���^c�>G�4���G�Tۨw������5��s���q��?��hLL5)W�9�м�N��2B�;��!K��v���LLaH�$�����;���]�/�J.u�Q������a���ǉ:�$�>��"`��ܳ��<L+�l`�u
�w���Dyߡ�}1 �S��A������'̤��;|n���g��"[ dF6���1쭡�C�u-��9��r����J�)s\k:�z�R�p����z�c�����m�֚Zh$ �P������KĊ���UYo�5�2��)B��[�ҸP���n���*o��hY�%��P^��
A_��	��J���
��-���V̵Ƹ��)��o�K#BG�c���?A�&j��)�<J�i���*QQ����Ek?��JH0����`f�X�
�4�4#�P�YyR��O*��hq�;@OIjV��k�
�@W�Wv�D��Ս���Y��a}Kc�(s�ˡ�{�i�?Z�y��%��*{z�E�9|��۶�Tu+��,�]�~��CH����9G�S1�˄��&�k=�$�A�@�DdB���"h��n>����%�XW�k�$Q{��٭��\�F��ϕ�V{�i�)P�MU�mP���vW`\Z�ý��.�b�����a:��H?�Ot�:�v�a���r�T����ov����{��V�g$~�Yr�a�J�,�/�B����yn��Ů	�l��y�KQ/��5f�?��t�������.�-��ⲯC����̹��6-T~���W���4�zQ�ʉ��I�ʠ�qf�7-�2h�p�a����q*�w��Fcv�JUS���v{��a����f��(�2��	s�?�cE>���R�4�$��o3
��n�o��l���n���	rt�ҙ����IP��L�*~i*�hCk��?yaq��{��<�{ZC�{*�2`�";?����id'��_Õ���g=��H\Ȼ�ɼu\���ă���&��P�ǀԏ��_,x��"���6�P:Wp+���L��g�'��g��ʝ sž�a�b�0m��fγ��+ �.8�d�k��Գ���z��̋��0n�7u۾�qR��q�{�<�6�İm=���x��?E��!!��6g�ws|F=M{qq�^��;�0�b�!t.�Ӏg_��zYKO;�#���K�ɦ4#�ͪ=�tJQy愊S���ľ4��H�H��c��郼�0V��'���AG��5B�4i!r�Tj�E��Q"3�"� 7	 &>���O���ɥ5��:q��Z|/A>���Ǣj6[��RiO�/��2,��tL����ˤ�)���DV�lQ�,��>?6�W�v~�"X����a������څ�A���PPr�m+G{'��.�LӉ���Ѥ�z�8�5��=%0�b_zy@�4lۭFi���
�{��ym�����¸/�4[�?�-T	�gX\�E.]�\� ��-*�=�h���۞)�"�՜���h��/�E��RǛ��Nɭ���G�,�*��E����~@uNf���+lKƼ���Ls��2�<�����/	:l��;^p�`��Pw�0�&����A@υ�E�"O �%��?�w������4)�J���ثg�t!F�v��!��G{�Q���s��fU�\ګ5�T����r���sA�RWE��>��S�|��85#��ڛ��/����{�2S�۪6U
�#�!�V�����`���0�4���+�wi��[���ɍ#�}�ɘ�)���zw�:Ѽ��'������.�ɌC��s�H�V��ʌ�L��F��j�?S�c/�QSR.�C�X=r:0���I1�w(��5�"��Y[��<��i��~�H��Mg��@]��K��t �B8hi�-��Ӡ�:�g�q�
h�n�w@����F�U>��0A]����ly���`����B��e�U>\iX8�DWz��o4lm�Մ�*��6����=1��L��Up�]|��6$LȸC���0g��z��74���TQ�ŚՇ!���{.��%KxO�\
X� ���=��;t�i��{�i3lq�lt?����Ŧ+]-����ɛ"_&��TU˯��j��W�<ΐB�U�P`	�gnUC,/�/�l���t�%��z���y�?��E�� ˕
���h�[�FE�J���S&�<�y7���-�>��Rp:��v�����R�;+<��h=���P������� pl��즼o���l{��;��?]������^�M����$pQ��-�!���~�/��?3}���ɆC-�^�aMĳ	2V�s� &W�I�wT�5�h�S�h�W�'A���G: �Ob ��,_�=?2^C���Tieq�%��}�WH�� �L;�)�-nF�Yb�Q�����˻g;�j�S�_cWSpz�ɴ�7'؏
�������P(�{�*����Q�R�?�FQ�9%v���q��,�{<������$r;��ר������M�O��|#�jk��`,n�-�u�$b��|������s��h�&3/&�1d�n�R͜�� "+�,���C�r2%DX3�$h�9�xk�?�d8�Kya�kcH���<�d��+hH��m��=�1!�����÷�s4�ȱ��+`[�Tj�K��2�1�T���id۽êl���Y�5_f:��t�����C-�^7�ec�b� �T�*�m!U%Ha]�� ��)��h�O�B�{�k,�cw\x�[�?R�6nQU�7���%�S}��%���P�w�房�d�	�����1I������[�Wg��BZ��PW!t��$f�wjx�d3p��ͭ�X�����v��������qT�����d��"e��$
�-���*>6�
}~Q���/��Gw#�4[�!�Ë̦E�equ�g$?6r	>���ö?�V����Bud��C��m����[HF�]�g�Ԫ�\B�aDf���qn�[�Lț�a�*
�r�,֗�0�f!zN!+�S5N�ݝI�c�@+�[�%��i�3}� ђq2:�'[�l���&
��HkX^�J�Vs3W�6��ݝE�n�d_V�^O(��J�C̢�g���n{��M⭜�\˕݈���_��	8���u-�G�Fgr��r�����w�_���Hg����9RpɇQ��T��ǂ��-�Q��
�ItWz�;��H�f=���5�\�<�-���s��5�P5!`r#]ٌ��,G3w�����g߇5�<0��"�,N�C^��7*?#���=W���w+�r����6���C��KPZ1��0w�M9��uy�H~S�y����qW?����U}���vwq$�[���r*�\�5!u�$����h*I�!%�8��B����#��(������Ƶ�2s��6�mۏ��2�'}g倈�-��e^��:(rjJD_���i�L7��:����њ��J}UR�+@g� t`���r&����1�&o	�{�r�95;cc=P�M�L8�Fq�o��:�����s��O��F�k��	]n����[���Oj��U.�r�f��2�IQ3�Xc��qQp��k��y�z��*r��é���߁p��V敜��,ޡp߀��������B҇�����%��L,v̉�n*���]�(;�H�ߡ��E��kS-�����d<:��8�H��7fk���� �ol�7`y�Pl�3�~,GA��+n?�+�v�4T^������}}��?�;���u��iKG5e����)���P�9	�$�#�>Ws��Xڴ\�N�q��˟��7��8��Uv�� �:��|D�X!�2F�Ј���Ted{���I��I�+�����_�ROS)�Y��f�����E'�5f���"��s�kB��M����Kd9L��%�R����J%�G'�|�:�m�+vzTJ��^�5��v��Vq��?�����e^�VC��H���ظ���'��n)��sR��+ѠAq�f>��S�fX�48$$�wQzV��bk�L[z�H�Ua�p��ʘy�D���@�jX;��!U���;(b�Q��G�8���Qm�����l:h�m�:å�"����?]�u�u,���?o�T�D ���xY��?%�^ifB���UC��ۃ��hC5�&x��_bM4d�s`D�ֺ�^u��QAy�FvQ���@���������z�Q9%�o��W4 ���}?�s���<�>s�~�qȢ��6'|=���T7�|�C��!R�O�\/�9���8?�LLa|bNv��}+E�*iZ�D�K�Q������惚�V�C�~ߞI]1/��.�j�jh^����U ����JR�B�]k'#�����&e����\�L��_°���IW��J2����7�]I\�PY���y�� ����D.�T���V���w-���e��|�p,��ʝ�@�P�?0Չ٠|e�F\M��Q޻h���7�nI�h%��\<��E���ڦ��ٿ|�&�5^e�˽������Z�綎�Ey^� e�����#&�UK*m+�|s��ȗ�=K��,�{�����������g�Z3�dԹo���.T�cKHLT����Ux1��v�2�<	�MB�A�4�����&
m��~��G�I�{�Gf�[ȸm$��m��a��ObPcҠ�f�e�G�Jv��|����ϸ��yU(d/�EP�����]�ͽ��eG*�`�
�?�w��b����%gJu��v?�Q˶5:G�x�)�,!����s���*��o
�۪s"{�&�8���Z]����]�(�����k�4���p?s�~ϛ������ӣi˻Z���2�!{��3�w������zqH�$pڪ�?-H���S���.+T�?�[�!��6���%���t���UB҇��Q5�U�M��6�9>zv�!��?,��83����{XL���?-Njg\��@�ǉk@rИ�_�@�\�Q��fe�Gb�`���պ*��Q����1�-1Š�.����~��e!&����ǳO��!6
p?T�	�.:q�BukpSO'�x{��#��4V^0��U|�d�E�}��Ѣ�,�ޫ4�Vb+�Q�l��Bx:g��b�J\�[�IN�#�������1_��ג��S��඘?���g`���Y{���&I���4԰��6��1F����D�uc����E$�~�vۊ��H`�AZ��!����aE��	c����� �3��ѿ�gUV�ݝ��� ���V �p�����S�fh��E/��x����TT!7��x�J+e?hӧ�)�s���i�q���+��!���m'�߄z<�����u!��Փ�Řߺs��[�?Ӎ��k��S���Ǡt���S"3��8UA����V#���{e�����uH�]�Q�[9M��f��]b|3�4�ɻ�<`82�Ja<-c��"A/��~�O���XZ/~��ԯ���N��iV��}16oD���s� ��v����e-��$�W�TV��=RvU�@V(�pD�	�����f���~^����٫<g�u��,.��ÄC��X�<�~��N<+��>���K��BV�Uk�[\1�_\�T�E-V�cǃ$!��(���"��;.?�I�U�~���i ���X�v	��� o�"���0F���^-e���������"���st��kr�2�8U�%ę"��V���V"MA��M+�},�2���9Y�}����۾� �1\vJ�Ɛv�}~���<���a����%�R�?�D0u��/�"�Q��6j��<��Vld�!?�I�S��ˡ��g�u~,�ot��x�+���4Xv�P�
��:����϶������ؐ�bio�f\����N��	�bz=��vu������}]` �\v#����9���V�(+G�����R��ܧ�^���~��]�,vy
��K�p`H�h�n�L�D
�&�Vt�����J����{�bE�ow8=H�T$����� ��Y��TJ>�8�J���C��ΰ�R���F�B�������XW��-@�d����	\�O�x/zLc���Z��Y�>:�|��B��H\2��[&E@�RB�5&�������� �<�'��
ZXGI�lk���rpZ��g!&o�_�#��op>4{C��^2�<��7�)F;��7�Ҵ#�W��3��8�.מ���:�vɞ�kDϯn�D���!�i���f��M���]��V��94��W��|�[��<�����ռ���V�l��_*�����p�BOF�P��w5�{3�օTCB�����*�����n+8R�(G�!i鐞v���d�Id�#М՗:e����ƀ!ǧ��;�$,�;��I���Z�FH�ZRu��=�<��,�uk X;Mx�՗�J-�:��#\�l�Rd^�^iA�M���y�D�0����m1�<�53�����lH��TƜY��NZ$��"�����j���e+����6 �����sr�wU6��짶������(#���?iK#���^X���D$�؄f����	 �Z�*uE
ܸ�eS[MQl9��h�V2:Gד�S��8:Ch E�u�c��/m�l�D�hif��f���[���S�j(�' C3�e�_GC>$���(���$-w�6N�c+��b�n�!�q�� ���Ɍ������^{oL�H4���M����I�b����q�)��J���s�IF�%��nG��9����>~��1��d�ڇ��xkź �wU[�'��{�ޤA��3�z[�tS�
|ͱ�{��>���nG���g�2?Zb�Q�-��
�`���,�&p�6p����d�J��1'h�g�4-H��aУo�#��,I8�K��G�Yj�	�~�9p1�%`q��E('�#���k�n}��S���.f8�FT��C1 z������}
���[?�"��k����er�D�g�XGa��0D ��6����ꋉ}j����$��ݒ4�'>�qpp��5�]L&sK�Ж�0aO�?�;fEi��������r�=�:͖Mp+��s؃y��J��8mm�"�J��j��KK�(�T��AU@�Vt��-_}M���;�]3P�b��M��w�X����V�5�B�_���z�V�aY�X��<�������$�P[��G���dQ�k� ��t��!����y�5���O��n�T���N��GG�g�j�y��*G<�k���vژ�b�!�iI�,WR�P���Q½4J�'�X���&]5�X ���줻��?�|
cey��qe
�`E�Q�+D����7�}._�����m~���砼�|�{ϥl��E����}���X~�@vW|�����T%�#Q�h�W�s��;�h��N����K�5�ܞ��`is�9��d� �(�{M��R7�qER`6��t;N��8׋!~�:U����#�+�'�qWi}���A#_@���>�J��>��2�Z�'fV��7'sW������H���V.e��R��ЫI�?[A�g��N0�!u�8��\���C�ZN|]��	b>&	'�Mn�HB.��i����ڸ��oB����"@rej��xӨ���x}W�D��U����..�%����|AqC��v~�ڡTʤ���{mj�
kc<n'�/
P>�+m�٧�I5�l�dYM?�e�N�}��/�������<�����`P�w��� K�m����n�eQ��n}CG��`C�2D3�����	��S�	��f�����L�al�ɮ�<[/��j��O�nq��t䞤|?�A���6�4i�nQd���x�{�U�N:bE��D�F9B7b�ű�s�4�ӟ�D;��x"T�-n�H��q�xq~���8+�~uKS+XkT���'O��K�#;��ʬ�Y���lzVT�q�8&�����AΏq��9+a�c#�hc��£�x���%*̙�%l���sJ�d(tT&��q�v��s�i*��y���
�W�e�IXY	�"�|�_�h:ZY��TK;fSDl;��pĬȰ����
��Cˈ����F�5^����� ��S�Itf�-Ȧ[��[��{$����O�+�!�=�2�ӟV�<~&7Fh�Nx�L3'h�!иo{G��11臒q�}V/�����~c::�b�mN�u�}���@�)��鋠��BR��s [DH�f+��~��4�ؒRe&�w�^je��|yV�&7���[�q�,e-ZiϏ�Z��O�4�,��=o ���u�y �d
2u�"Qm�+��Iq�C�%�ڈ9��dRh΄����ƕ7�c���t����eiܖ2&����n�D��T5����ˎ3|G�o엥1P����h_3�˥���,�wIr�PA�ݑ,�;���;��%�hw�ψ0�ҳ�&�S�X��v�@��9����,ξr]�<՚��i�� A�a��x���vjš`6���)�<eK�N� �*B�Ђ��%UH_���u	!��h�m��~�)�y:��U�%p��=�)������݊r�,��X\�C�-{[A�]�?
��e��6�z�nU*�8=�9���,}����WM<��4�xkPt�a�E��]��1�/L��K'���q�[��;q02���^T?�ĨZ��.�9�~��3�����ZE�&�}��U�=_42������Rá�����&�f�b��۹�*m�}X�$� �	��.���H>u�F1Řx'�{'�p���^��*뜊)��Dhd-�]>"G��
(L�����T�ִ�ꄱsb��r���q��k��]�aw�g_9|���f�i�H\k�.F��2T�u�k�R��3��+KCMf�Q[ml���*Þ8靳�����˘��S�A~��h�)|���_��5<[Ս���j 2c���t�����[t�rɄ�"�5����E����8)saA��bK�#�oy��x/���MBݺ=����@%{x��~u���bO
[��R���y��$C,�-�G씩c�JQ�m"0�!�d�/9��#��f��ŗ���>�?����ѷ0Փm�"@P�b�M{�LY���̪��En.��XW�	$�تc�M\�[`����{28d��^xe�!9-J7>~��w��U�8��`��I�x�#��~��w���36F���"
�C��7UѮ^�d�[�5*u�	Z%'f�|����C��+��LEF��,�^��Zj�u=���א�4dĽy��b��gB�LA@3rGsl�%���� U]���_��T���u��B��:�rA���ٛ���}�^��%/}f�\ 4��S%�@Kw�z+��M2�'��FG�Kr��;�S�
�S�v��/v;zpH��
LO��1o���
��
)̾�c�1E�ڭuB9@�}q�e���S�]7���A%D�l�D�:%N�\Dq�,���ݘ
^��)�"�Q��#����u\���d�D��x{ڐ{]��rG�S���>�M��7s�%�n!�<�ZM��&Qx� �6��?�lW-�J<`\D���KZ��h��P� E��h��Vt�g��ʩ��Tg�� Z�0��z�ܪg����f�(1Q��7�G��nWkT�g�M�Exkҹ�??;�j���m�����X��.�m�W���;��Z(HN@oz��O�.�Iy�=\Ѡ.���p���na�y��<4믌�8�&E@w�1�v�W�e�"�϶�v㓊Y�Z��J:���LdY�R��V�<�+'grw&&��R!Vl%4gzG�no~v��(���*�h��L]'Tq8���v�������N~�i����#H ѩ�6 ��P1c����D�EyJ�#jdh/�3��O�X������8�PCu���d��)�P��	�-!؜�C[�J5*������r���������<5	�{̭���$l�YbL�̏���ւQP��i���e���l�Z(�|�ăv�����*�9���Ѳ�S��6�wD��^����.�J���#W��î	26�K�C�����ʃw����-��<���}���Q��c���Xfx�"65����F��-�2Y��q��e���r;Lp����k�@�55�}��(po~�z��l�Zoc�͜]��H�Qra|et� ��w=�����kD�����]~G�j�^b��̮YƔ���'��M �Vu����5��i�
�+N�~��j�r�����t݃� �)	��55��>��)����4�Oɗ��Ͱ��[�uF�D��W��t�+�2�\�<oЪ��r��T,i��P2��`�A�DX5ߜSh�b���2��q���$��I�LJ�L!��6I����o4Sm�9�y �A�<�C]�CY����q�"�Q�y^�6�뤷� �RN�r�����%dL;O�s���
�9Q!?l�\'�	�S�M^�LQ�\G��C�G]����V��=miH��m��BĠ�M���\��$ �p��;�;��\�d�D�����)u^:!7����d+)/�:�Y�J�%H��}%��̈$��e�@�ʝ�nE0[ƽ��؈4���f7�NȲ���*�P��"ҴVI��'��}�ĿY�`�=F���gު��B%�����+Z��ׅ�݈z�j6�T+r%�q
_���ނ���_�?�sc���3O��\�r?�l�#=iT(�!�f�5[�e��+5\.�q�%�J;�o�yl�q��i�]\��
���+�,>�^^�ٗQ�@�k���߈�k��㜎?�#����i�j�^�iޛ�h�:B�5@W��6��9�Byho��*mWj��[�O�!��hf,��%n��os��>�����r׽���^��7�F���0�y���@�/ޓ�@��ϒ�Ğu��U�D�!�t���a���2s#b�����w�΍��Xܰ�ɷ<�4*��-����� W@�� G��"�
1�O` 1�ѥ��be��/��Ee��a��Uj^�X����M	��`N=���@�M$�XL=M$b	� 0��|�g��\M��q9<3_��1����@ꭿ��a��(�A>f���|�7��W�%:���r'Gq �"���BR|I�<	V3ìZ>�[�67�t?��������\$'@�;2�oVǯ����EMYiY����2���+���p�"ݠfqb���+6R�OG���처���.�I=���d�`�hܾ�ɨm|���ьʻؗ���V��&:��	CW%J�u��	�pt��*U���	5I��uq�4k��E�R�919l�#�'���IE�f��?��7�	�ea�[�����Gks~ z��]x�n_�{��q��wR+��B���ѥ�b�6_<Y�}ڊ"̷�Zr;/r�s�Һ��HZy)�u�]���g�: ����Jf�O}�}�.��r�CGU��F\��~)����C���|���A:n/��0�_�9AE}�V��8���%�Y�P Dc�����}���
�I ����Ԇ�+������픺7G,��oh��\
J�M��[��Ki�?�.�z��) 4C�P��OzڅF<
��dt��FECP�g�w���C[h�!�����#T�tH F���^��8��1^�������17���r��X�x�&��H�N�Qi~v���CuQ2Z�]-h��V���Tg������Ď��uz��/ƪ[HC}�xzdgp'����,6�V[X��g�r�%tj�(o�ǷvPe���[�yTZW7�ǝ�����D	Q��ZY(w�L�:�n�z+�5ށ��R�V2�\�(�:{q�G��G�ln-�rt�8^A�#���c`��L6�l#=���p�9��d���0Z%	1G�P>��U��h�L��N��y���^�7��Wg����r+����|X�������k�<�_�yZ���]����_9�?��]�_����1x*���GPE�羑�۟]Js��̬��/���bM��F��U-J�����
�a^�Q��7`ip�Zs��ڹNUka�E��!w|��.69� ?�OAM��)e i�p@h�ٛ<I�d|�,WLm�5�z��:��x ��!�{�W�}���8{(�@����k��#�Y��]�/�����	U��|�<v�M���s,C�/ܢ�\5"Ql��9�2i9qGZ5,G��~`^��P���V���
z|͌,`Fe�%�{�ioI?�~Q��z ����N���PF�.? �����,O��mT/`�N� Nu��h��N�{�-m4�rB�~��".L��#���`�p���-_��� J7������<ޛ�>���u����r� �*va�b7Z�;���֌�=�R\���qߚ�&��LQ�y���l\)?Qٚ�ވ�щ��q΁ȉ0�(����&�T���F���E��眹��-꘥!�}�:7��(Q���t��U6X��U�ԛ��{�Y���
<��l�;1�oy_�������f};�1�����x������8�ɧ�N�^�Q"1���Lҹ��}9��0!J�qz-�D��O{����=�%M�{�V. ��j)k5�e����-�+��{�1ƄhZC[C���h�2�9��D&��C.Eq7d�F��%$�D�O�Yc�a��E���=�9����*$	�7�_9�9�}��-��i�l��c�tKg��1m%�Z��.������������O���	N�h;�R<E���.���(�K��R5ȦZ�Xߜ�l9|G�Yj/R78�k��hN��cO��p�����Q�7
J�P�鸙z~�?��AΈ��t�T�H�&-=���.��,8�k��W���ͨ��6�4��A[�(<�������?�KE54o����3hd� Gy.��)׫��¨�d� ��֮D���aM��c���K��`���m��1 _>b�%��s����y��cd��MӤ��y���b�����>��iPw���Pi��a|��I|�`P�L�>@S��	�q2�.&���;:�"&5�#n�ڠ�N8��[I3��j$��<�y�7ɩ)���ӊ��u�q$� �i+�'���tMjs.}S ��2 �j�V���C������O�����.��g�/�Oð$g��V�C�~�����Mŵ*"~�L�r�w��'
�7����uyvK��?�_��YT��Y�_RG���;K��ng7+��Iw�2GKuH��Um��>�g縴�G[�#Jy>�Bc-�(q�ރH>�T-R4���� �GJL����]s619	�R�A��Ƨi̝r3P7��b�R�yc��ɮ_�N��	��4~���HP���Y9�&�پ�^�f��0��߸;��pYM��N��:����Ub[Z,ǝ;��K��,Q���s�W�H$j�=��gv�xѫ;�Id�0��m��ӵ.K��v�z�E�9��ON��voG�-N�ii�Ʈ�rR�6E%u-2��T��D�埴۸d��t�����K�j%YX��l!_>���j�g�.\���f�6mF��b�_ԛ$vE���l���������W���ȷg$������sJݶ���|�3B�O/�\��U���w����W�1_bMځw����Q�B����Q6��A��P���z����ل�*��1�@tY��:i��4PbRCI�Py 1��NS�b�9ݔ�f5�e��8м��<�"kd����Ȕ�_<(;���:� MGhu1�{"�Ԝ�3u����AQ��O nv�V�Ie��[jq�5�^}���������
px��N� �P(�=H��ۘȍ���}4����4�:=kA��>n��d�8�4�{�j��'Xx�cFm˽���Sc$?�%FO�kD�/؍ݩ�WC]*A'�#�#�@�_j_��G��UB�/�Q�4�J�#]U}T,)y�k�:G�R4��?�jD�\��\'����+`��G��1+���<i�ܵ<��ؤ4,��1��K8��Y�̨��Q�M1O@�G���`M�U���w�ءB�rR.�����+
z'^7�E�}�� �Q�@�[o��i�$��t�T?"���z��4	�	��-�$����� 7Gя���1��J�@�v��8�ͤz5k�8�d��"u7d3��\!]SN~B9Gn��Pm�-��n�+
���d��!�yKYM�e�҈SF�tzf��LM*!��2���=��p}83��ό����mL�b�S�O7����Ѿ0ص�ѥ�ܸ�+�H�}ȱ��x�$��[!��5��	@�f: �#UDz��r�����bW���~2����Wdo/i�tȊ�\e��'Ă*p:{�+5��Q��9p�\���N`��m�e��ݍ��K6���R�,�e�ŜB�>w�GH��C<	���1Y��aG)�Lc��q�GUY^�nU�B
9ύ����{��~Nӝ?���� c��'S�Lt{2K��Ɍ�-@�-��Y�-��ӎ�������3����lSfq�� �O%���2�5_�3������;�?B�ί�I�
*�	���~h�<$���x��S�fι�yґ���UD�I���s y�z�G����7�}k��[=�$p8?�g��5c`����Go7���҅�~�� �TZ�5u�8Eb̽-�L�����}|��9���kK�ݼ&��M�flMLK�;_9Iq�M�����5��<��P�C�a�E��n��c�ɲ�G]�J�E�"8��),z�0��p�̨e�x�����l�
��t8����
�r($p\'\6�8�d����ea
No�ܼ+uɈ�^�s�.��U,3��ٮcm�EyŚ���x0� ����L g�{�3��o"� :��B��׃Ŏ�vxp�[ �FU���p�*I��[�4�%G��;"4�O!_�%�^A[.ٿ�z��l��1�j�	��RzM얁���щ+���J?��ó�y�h��2��o�B��8ꕕ`��D�WN��Wi>B�c8}�bY���!�rY���o��L�+�N��*o��u����F�RJ�����-��h|v�܎�p��%to<D+���4A���G=R�+�p�S���J�k�rxV"*	�L�{Z��Sw�'���]�<�)IĤ��jy7���A_��T�����o���Jʪ@u��޸w/1\-��C�r��IW��O7,]ه�*���d���!�{��>���,�Xޣ�A8�|L��R�0"�B�~#����?�&�]�![i���K������B<N?%P6fߘ���C)�n����;c~GG�zw����P�v3u�/v{�!��F1��k]���N�Ҵ����b�����7�)ɀ|�������e%ͭ	caJ�]���w����-�#�����٤:��o,^X����O��9�޶���J����c��v�@��[�dż����׼u���V>/6@�>�4�;����g���.���~�����4Z�0�*�*0`�1p&������ʘe������W�b��h�!u?}#G����0u���T�s�&�G�Y�|�	��	���m�.\��k6�퍏�o��`���w&���2�l������Rc��`�mI���
�v�Gb�,�b���#Lsv�G�DC%ƽ���ĵ�?Ҥ6ig��bgi�R������O�!\V�P��A�IU���9ֹ��1:��.�`�����:G�7x����;P��/.F�!�%?��A
�A���j�|��sW�`Zx����q��\�~���s�� ֛�.�=[�`�	�p�6;��߱I�� �})�+��LM�S�V�^�0j�oӆ��U�6j����Tk��s<���c�4I6��3LCy+��x����|_L�����Q��^}��*�� љ<�Aho�~�E6j=� �t"��uJB�O�)-1=#�g�� �?H��aCӞ���m[�E:����:��OΫCm� �R t.��U,��m S��ˮ;(��VC���eK���L�A��{,ߓ~8�}&�'?-��5_,%[ķ\��2��A;�����o�u����s����=.���&~w���lй�TӂrI�k+c�
"w��D=���E����ۤ�,�~�ɴ�u�a�L/�	���u��%+g��3���;�V��k����KU¡U�G�mO~�f��wO�o%�:&��N��������je�������b)��*.�w_X
*����̪��1��3��<$g���k��
�o�$SS�
>-a&��
0�+����$�]��=�F�&��x��!naM�kB���Edo�%�q5����@C�Qw���B�{�4���Gfu�!"�R��Sd9l���Q�Xm3�
�Tq���hof�W��,�RX�ݕő�� ��`�X�ð݉N>�\/ ��D���l50����:�z&߅__����=%f���S��P�����g�5�������;|l��P���H����ꮇs�\ɤ��o�.�
�\`B��o>����؎fH��m�.���e���0[pz�A�=n���+�8�\5���%ˑ���^��D\s����g(/�L
�0�Zw����S{X��G�����H�zcv�U�oF�|Cl�>py��r��^?;?97��+�:^����%B"�J,�y�q�C4�}Ɏ^Q�fqf�����IGd�-p����o��C���L;� ޭ���T���L�J��Io�H�p���/�b6��8���f�l��d�ɹT�WA���}SL��;ݯ��c���.��Qv&�w��y�b�R2#lH�퍅oZx~&�C�L]��J�~�����H'���J�J1L�7�Qw�������5��D\����?��'?W!J\���I����C�<�d�K9�7X`�9$"�B|(T ۓ��B�Pԥ	��c8q�d�1͵�fl��r��Ũ�u�[>��`i��)f�����`�1`�pL��>׺�[�B7���Z͗X�Wb.Gֶk�FCh烃���Z�2�6��B�0P��*Me�4-t�ǘ��1��]6� ��B[c`m��v�rZ���ҰF_4o�G[<��e��VRj��`�������݉>�?�J;�.��ce�_
r�@��s�Cs�Z��+=�_m������[�$u�$��ϝQ�/[N[ox�&���9E�U�	0�;�,��+x}�`X�G<4biw���9���Q�|�Ub���p�t# �6�&)Z�U���<6c���]FCq�r*�K:������S�q�`����a�y����G����)������T́�j�9.��)�bO-�/V��Ԝ��PX �ٽ�D��9�Z�-�x��GG �Z�o�x�F���1W]?��;��X%J�~�3��w�R�,�~�>�Y��ϐOb��.^��L�U%����/�N�>��6]�:���P��l	�2�Պ0�Gu��s��Z
��+Ԏ�Lʎ��'h��y��L�V&"0�K{�!�v�������Z�S�.q���	3�I)w������MZ��1FZ��≏ޛd��I�aX���M��9��&��|x�^o-t�张�)i�v�7|�� !8� 2�a//�4Տ8�'�w��鸨�o�1��e����z&�@�~�4���
��L����}��&,tu�ku49��,3��Rl��Z�e��sLՃ�F>�D�4XC�헟����3���	<��{�p��y�۝�L�5��Dfm'��%���{
���gpb7,U� H~�����n`
E�yg�7oK29V�p�0�f��Q1R�G��w@q�EoECn�XsA����~��O8Ժ8l�����
&�B�>�XU�&�9*��Z�/Z=G���Ȭ#�d蠊3 =y�\?��E��ک-s%��U��>��!,�9 ��]x�	���e�
ĤR�j_�D����;w� �Nh����Oޠ[O�(��ډ*���%�=4@����l�
\XW�`��$�$�Z4��L�x�&T��
w�f�&�%$��s�����`^�u3�"?������uU_Ǩ �T�%�r"PV��ޕ�Y4�����6&
�A7Έ]3�Y x�[ �:�>xE-S*`�'	��I��~Ǆ���!� .��1\k�rGCDm �7}��JD������t̀�)��@�bK��	0_�z��\@��b��&�$c��BO�@}J7�1R�Z|� �!�h1u��S%4￿0fa�BI�@i�+Eh�!K�����K*�c�N��z|�j��6hbd6�ɤ9�m�W�p�>6�fW� *Y��#u��9�`�R�wE�3 �0ĿN+�~qlc!}cy��[Xͦ����HP��D��Ml}	6���ܺ�K���&=Q��̑�:2���C�=o?pPv!�-<��Y�����c�o]J��S�M8z�7ʲARId���R�)Ɖ�,=����`��-�����u�6%�e���j��ʃ�ݧu��$��$�M�� ��3�߷cI2npHғΛ`殆�����*�s���V���\/4$����p-H�&b��z��6	ާ��4�<MR�Ўø9�ʥ�2kO$04�A­Q�&���Dm��E�Ĭy��$��kvk�pA����k����$U+�6?;�CY]?�ۜ���=��0� k�,�� F��(��o�Irl�Dܳ�e�ϫ�9��[v�k�Pʀe�����0�oF�1X�d�컩?���0�aɂ.��/�
����$}Fte�Rj�莶������
�Dt���=�x�~� �x�����3��J �E<�x�ndN΋��&*N^b4��3h(���ĸ�y |�b_UilpvK���;��[�������{�H����}\���"f�z���&�J=��H��L�����!r�q�zُ��Ƈݮ��"���M�@�������{w� L}i3�12�(u�e��d�"_@"��.�n~)2�yI�>B���l�Jg61��h��e{���!�����1E��,�|�V�'�Ԗ2ۜط�;oB-k���Ѻ:��a5|��$;��Z�>JԄ8��o ������>�T⩃�3���ř8��>�7�`�]�R�˄;�ۻy�S��^|;^�aW�r�j��03�N꫌
UۓX�r��&�Y�_ʵ
�p�r+5��ܲ(�?�����o1@����i%�59 {��#�3+*��}����t?׆N��'����X��a4�Ev��vے��'S�%D&�{|uh�]\(������o��l.L�ج�Z_J?�j����A���z"��l
�潋�Y[�����f]w�W�"9����}J|2�̬��)�>�낳6���@�t�=�r}]Ul�4���l�P0m)�<�4I8x'�-����M/���)m��C�4ȸ�W�V���{s��4�����̔�yb�֦܊�{��1�h��UHN	��ڤ���mJ:D.x�4����y�Đ�Z�e����BuPj��g��@���?i����*_2D$��k��	��*DLcQ��<20����{>���l�'?=�+_�Ȉ�t�.�*�&�}�{��/)��d�G�s{��3/kG�{T��/�***MY�|���s 3�e�E��<����.t"�=8�O'	@�h9 ��,1kRm�j�?��r���Ǩ�ϲ�_3��T�HO��օF�|�٢	н�Sө���Ew�ZL����᫝�jL��0�i6��6�#�c�`�6�V�QGE;<1K����ƛ$���=�����b��;�^#�&�b�*�w�����cKT�t�C��N�OA��C���v�P7ꌬ����0g�X���Mx�m&�.��鏣h?���"�ka%6v}V��yl��	GdJ�=O͗�?-' �ڢ�&��N�V�.��l&{��37Jca����.�<����g�dٕ��d���5���7���
1�IOŚ#�g���:�{��&��L��:A����y����^�$�0"��+��p��9�Aɹ�����Y��|%��R���qؚ�t�����F�!��&�Ǻ��`��Zq����D�5�d�cC�+�������I�e��LE;��Pߔ[l�vPJ�� �Z�z>B��J��F؉��&s;W�Y���]Q2�Ҳ�a^H��iak��W���"�[�a��jb�/�-@ /��$�ܢ���z�����?��5|����{]Y���?q�R��=������	�ߍ��#�|�㎏�� m�w���D�t��V���$��څW��(79��@1�6ZBK����|>���ȏ�������S3[ OҦ�g`���vH���B�ܸ����^2tFc$����l��>�9�k��Q�#��V,�YL#�����xJ��d�?�ډ=E��M�9@�=BO�F_���飩!K��'�:���h5��_��;"+ha�S&m��Y%'J�h�0.:�����_�G����"ީ���Hv'��(��Z�j]�5v�2��5,�@\/��y�F*H�Jn��GC-:!��{�V6L�DxO�%5�X	K9�}c�������j��w֯���rx�{@�Eк���=�ۚ��@*�S� �6�ݍ���2�X�s�dpA��!�m�����(:x�ϋS1��\�R��%��4#l�-�90L5 ���Z���%5)��
3�-%Ѡ��0
,�_��+�3k���lI��)�@d��z�Zi�g��㔆�-�!����7�bUIyU�n�*bЍ"(6�X#&�6BHː�E	\�t�x�	9�@o25(U�^�w���š���{=4��I��D�\;'�"�䶰E���]�'�h^�$� F�	�,PL�*ahoM��b�<r�#.F:��~�©{fd��.�P���C4^�K��G���-"jv���cZ��wMi� ��K�80���e�,E��%!�+s��;!z{)#c��.^�[�4�S��wA�@����C%�'�
�}��?�M-+I��d�2�)#��?A�h
�^������+�hS=���"�����q�|cF����Ɂ��[�n@���/īG�F^Mw�j�jra��&:;�צ��MPC�.�-f0����A� mL�x��-A0�0̖�r���d�9� ���zOEm ��&��K�&[�E�c���vϭ���,)�lDC��}�����sQ���2T>)�X��F���Zۄ���U�`��NHS[�5GOGJ"3�j��*��A%����bO� +i��fc�CP]�O)�PӅ�ɉ*d�\���N����Gۢs@P˚w4���e�ޓ�'9�6�5d*�+��$���R&ZGR�ס�7�h�ힱy��d!�h0���W�J��B�v�6O���U�Yܑ|տ���?�T�c�f�  #B�� 4S ˱���r��]Ub@�ׇ�-b�fBJ^RT�ZM9�(+��p
Y�T&�F#��(&�w<���-��"�<'S'���6��j��{R�ʳX�y#�g��ci�NڋIv�T ������E��e�v 1K��;�롮���Bu���/�|?�:��,���叼'!��*�&%
�v4����o��$��3�mSH���0ϳ���+#8�'����95ԄyKBM�10Bҟ�3��-��z<֪� oM7w�>��l��X�nu�7�\E�s�D+2a=��G<+ٟ�Yk� �Suj�qHU�W89Z�������y���� �8y���
3����s�>�ŷ��U����޷gı������/J�ׯ0^͜�%���I|۝|s�H��5XC��!=��g�����_w���j�Y&����Vv�IabǛ�.'�,>ks��J`�ž�-�R�V�Y_L!�7�,��4Y;I��ֻ\���z
�A��l���k�LR��@��F� ���.�/d���nK��~��*i���wQDT��*,���csjIt2տԽAկ|��N�lf��E�����-�7��u�|ث�w�|E����E�Ú�#��z�4�X�ysZɄ�tT�+���%�n��5n�	Nax�vG�(�4Y����k�TO����Í�6\\П��l���H���!ǖ������ڧF�jb."�(9,4�:����KFC�����:��������ұ�VK?^��Ńg�_Vn�鿶
��f(�4�	^�3M �'�4�W��P�hĮ��xk����� �K�������{x6H�y��bS}�_�mKi-��I��B��J��N%���Y��)��S�_HQH��81��>o�\����y
����x$������1iQ���Ae2 F�	'&
XY�Y9ǊY���w�V	:��|G�x6��GW�S��b�L`��/i;��:}$�����3xc���B�h��Ż�g �fj! �!;��M�~Cw��y%��d�m^��2�J�$�_uy� σ��ή�%�s��-ٰ��l��ߥg��g�f����a%YzuF�kIqZ@o�]�_ɔ}��j��C	M9��cn�g/�ƪ��yF��Z�Giݼ�1��.�U֚-b�H�����j��*r��@p�/�O��k�[[FZ��i�����y<g-��B�&��[	L[;E��q=���"@HL�^E|�[��?��z �%���O���q14G�3�A&�g��1��W�!e���=���j��}�*\@�JG�U�>k���ƄU8b:���o�M���%R���0��GC��m��9^^M�S0$�F�+���5�601-E\�2�D(1ܚc��q�nb5��0��� �/�¸c���Z3A!�I�I�X��E���>�c���1�"�d�t���i�$�m��5G�
܁b�Yu�G�Jqq�ږ�]%ݪ�Sy�0X���)��!.�R�D	@@ɝ֢��:A�s����=���5�)��Խ�}��<&R-gf�`�,����o��o�.��9��59�J�I=ƨ&2� L�;A"~��(��-<Q@��?�Yq��A���$W�J�9R x�)�&��4�ڜ��.S��χZ�|��aU���]U��OǤ qOo�cM"��J� |��@\���N'S��^]�DiN�=�~'�����i�µ ;hm�Y�=�Cg���F������?6<7Ef�.�R�B(2�q��U�^3=��H�Ү����lI��X@8.B*^8"�Sd��[����w�@����:'Gw[+���o F�����P��1���o6ru߶��#���\�>Z����Ì��y���� $�=CF�`�F�җ�Tx¥3��.��5�o�.��JݐeF�P�禸Կv&x�9J����>��c�5jޯ�S�� �q*���s}�0�z;�oDl��/���:n�1{��&^o��>��`�����.',�c���%�f��w��� �om��HC��$��h��|R-��=�6�\���	�D�[1N�����b�{E�Z"��2t�/4���p=U��u4v3� -������B-�W�`9tQf�#�Pi�o��j�B������{Y?{����k� {}v'����I�-K��SO�X^3^W�v�����N�"}r�t��T.��!m}'�*���ſ�0mG�/��f��N�D^ !��˽x���ZeUR���� �~�@�Z�	3�/��탭����x�m��N�{�R������=��MM�Y�!l�6�^�J�XFF�'}|�B|�c[E��;����"��9e�3!�h�ʊ��B�|A�LL��F���;��$�Φ�F���HgVb����l�ϝ+����
�Y�0�%&����a4nة&;:ڥ�j�l����kj%���'�2�$|�n�;^ӜO�ᙀ4c=�⦮ ���mK~�|��hw_Y�����;�4�3��T����}����!��n1�՚�\������R��:o<��P�>!06�5���ks& W�b��Wzޮ���ĂЯ�t��C<�W7��o.)�����Y1���&w�e�[�� 42R�F��<���0��t$����V��t����Y��GY_aR�̙#�<OX	��C��ܣ��I�e��ڹ���QR���=)��,΄^�sh�{��}xc�k��r�`J�����pjn�Ƌl}u���S=��c�fWר�nk<����;����6�|��Xe�m?r�{�b�J�`M���v1î�"��%a��%��m~Er|�U�M82�设v�CJ��w^ �����Ӌ���|��/��.������Aq	x���Ժ�T7%�@c5�]^B��qеz���u �,��ZE��FmM
s�q��rb�d�(߇�H�X�*��0߾\N�[�K���AJ�T%]����;���>Äî��uN��CQœ���/F�-|��h�頻@ƒL?���)�kH,NGbfh� Õwu���Lz�r�c�UǍ(kW�V�8���P�s����Խ�g]y�.�}s��m4� J����09n�J���X�}�#����h��q�&.�!��g_�P?�y>B��h�/pF>�Ʈ�F/$D� ���KU��!Y��X?���j�G~��ق�&o�7\��&�`s�p�X���w_�]�|nCS���1����8@ Ċ�}Z1P�ܪK�`CEZ�BV�8��l����5I�me����� ��I��Ј�8(�j�_�: �D�e�V/[�b$�L䁵�=�FY�;U���@�r{�������sD_>���L�eq�$7�FS��G�
זV�2�n�va��3ߛ�Ȑ�$�<�{j����`��� ]���7��5���u�I�88��j�2��[���#c���,�w6�b��e�=���qL����nW��(�UKQ�Qۓ��t�n��i��Sg.���~B��"���&�D+�+�j�amX��''�X�����&�� ��3�����M��,A�՟*cN�p��h0B�`�Mf�>�!�m$�j>/����Q�-�[�WKЖ�pP���p{7٢i(bκ{c�n��$�h�AE!Y���I�=��Q�yWV��UpN�ꫭ/��'FutRQz��R}&�p۽��� <?���o�J�E�}4�����,���LKo$��&����쪆Xk�IcXG^FE�Rq��`�|���6C@U��Kݞ��Y��۰�����Ұ*��,��~o�/�%��l���F��g��x�T���v�#E�)�$M@��z��a��a%+ta�w3q���H@��x�b��O�O��V���'I��������7����+W�׸�:{�[���Q��w��+�����e����w#���2�ᏖZ�װP���d4�@}*+2�~r�![p؊Qp�SL :s(�.z������փ��yIG7��xOް}�/��	i��^÷��Tq�i+�Cv��P����zX��gK�'�5 �v��G?�o
y�K^CG�t ��n@�	�\xS�TT�#�ЧJ��r����/���t���.�#���pƍ�����b�\Q�'��W�8��|���� z��)N��IUJq�/,�(G��{��5ߎ�/��x�~���v�����ƷT��8G���B�fr�,�2�.�Me�Є�-�ŋ�u�ꋠ��㺁vW�sI�ĄɅ>]�z��܉Pd�+h�`H4��ir�P��0w��_ۂ1bӂ�����Γ1�L�w ����T<3t��|�_���c$�"Y���u�'��K�����[�V�b�`O^�t鬀�c��P���)��{�T4nM�1jF3��<!�O�|�"Kak��~
`:\��R��[#y�&8t���G�IӪ��*�����p����t���CZ���t���+J��,Vx;"e'��9s��d��	鎟�-3��L<٦$J�g�cԘh��� ?L��5ι,�2�#�f�{?`�r,��	�����0a��Go�Ɩ���Kw�l?E�V�0-��g-[~*����A!�^ϧ|y�́l� ���{C�c������PQ����?U� �J>��Zf�]��p��� ��x�%Kh�-��HU���qs9��g��~���9^6��?�q��2/E�<`	��7���j�����4��*���So�$WPw�ܬ��t>_"bd�mY��p��U����'�<��g�5ӓ�j�:���u7\��+�B�؁\�O2��t��0��]�@Wϸ��s��x6�K�B�J�����{�\b��g!��o" ��\�@�Q�,�9�o.Q����^� mZt�{X�у��rkKѪd�v�V椣�W��z��^�;>�0�I%G4=�K֓s\��V����I��p�ލ�v�3�q�z7���0&��`	��rhA5~��9��S�!������|_2e�\e4�z������Z�)N��%��ݭ/j%��⹞]"�	��c�.�.�X�L 	�N,�SR��	��đ��$�0��G9�A/O茴��DO����w΁�K�H�6�z�nu�K����ߕ�o7����繠�� vո���{FkM���k��z]rh���´z�dā�_���J0'�˰ԍ�Y��ӌ����xF0�1q�XPf� 6
���
8T~OF�0��CRY=,��}9��4ߡ.�_�����z
࠶����Se�V�N{��3cN�c)a}O�)�Ͻ��K�	Q,(.�A����D�WUg��(�;(���͙��|�x�,�r�< �P���ø��j�#W&䡪����eX�ܫ�z�$�Ʌ_Ph^
q�~h?�O,nܴ5N�~B"���e�>��Ni_2�m��~"ʞoOLъ��+f{G���T_m�Ҥ�U���F��>s�v������M� Y��cJd}˙z���K����U�2���H}D�9�5q&��l'`ֱ!�
�؉V�^Ѽ�k�[�3�u�z�l�P4륍�>/j����������Dcxӕ�@{�Xi��~�� � ���ދ�k�D��}`a���% ����7p߂	�� ����9<g.?JW1��C6
f���6��!��6̪�O�q���@�"��j%ƚz�G	�N�}ïg�A̭��";�w���	�i����vQ#�mD�B����9�Q�ӝ�w�+�wK��"d�x������U���[N���`&7
1#�K�5���206D:算c�r66^����_�@u������|Zu�3�����e} ^�;㊼�Q ��%�ƳIҔ[T��c)1����#�{)w���X�`M��J�>*�p�q]2)��{4צ��A�|#�r��]罕��J-qHf��C]r���tXwi-\?�^F�G�̇Zx��E�&'�Ev���f�D��F���C1%��\�y�*�M��\�-R>��X�������c�pK����X������Uw�R嶿��W��e��f"PC�B��I���Nw�7q������B}v�\1��,\?�"��Ј�1���*��k]�#�q!v�J	L�E}�6}]g�=|fQ�(�Mxs�Mm�l������3�y��}z�e����k/���m��z#RO�Iz�`L�;�S��:�n(u+��:T\�K�C��.{d�΀A�����v�;��@ʐ;?��M��R�}h�يR,��P:�~M;Yj~z�dBٹNʮS�3�N�G�޲���d�_8���'wi�i"�;��a�*��n7�cpA��^F�#T%��O��Ι�*<(Kz,zbd��kO�@پ8s�VDy�Ў[�w�QP�����Q��N,?�f=�׃�A]z�
� {"���D����m����0#�0�s4zW��`�������A&�_��:�#N}�	�8�VA[$��bm�+�:H�����.��%)�������r�b�Z�j�S��\� ��+E�V��A{:���}����z��=ќ
&�'D�8r ��cg����F��+�ь�a��4�qo뾪O@���\~Ķ��[O��%�!�1��@m�ݞz� h�g�Iݡ�f~أ���{�Q��$��G;�H��5TvǛhz���S��ۧ3G�\m%^�d�C�rU^�}ؿٲx K6eB��-/\n4�h�n*�aF ��慠�(�KB���5�EU_ܶ�ŅG1�"��C��V��l"�q���Q��N)�wa�M�N\OB�kd�D��_GS�t��
�K"
�U��J1g����NZ��L���E�d�~�����K��S�)�Bs�R˫�؜y����߃)�f������jH�ڒx�6��9`����=A��jz?�d��@����I@d��Vc�Q���=?tf��rG�v��de�J[�bb	q�K�:m��c�f�p巗G��~�,c�A0�~�'�A����π�����+!�g�΅�=��|A����� �V��m�0&���CNl^x�_�AQ#���D���Ȓ�\d��Y��Bl?O����Z�N���Ze%���
fV��Q���<�J3��ڿ��>d.煦t��L[D�[܈���(#"���`8�@��%�Jj�b�����*%�z�1���MA�׽|8I$�j%rf�+_��z��7�S���Q�ܱ�>��.o嚟x?/m��v�A��' ����<��%�h^�(��Y�\���0��U���6�11��:5�4�CAI<����.JO8� ��,ߏ�Y��D�����U��|�9�6cC�Ϛ�0p�*i+ͳ-A?��kMD���X+�ܧ�t�w���)��+Vk�W>\��&0\Z)e���QL�9��X���!�1o�%��a��v�Z��W�`|ձ�$+��e�spdi���ư�����b{+�)��%��ũ�"J���!�0Q��SX��>�c�����\��e�BgGa���iH�I�Nnã���]D��z�u؁v�:`�'��V���-���kC��8���l'L�I��7Z������(PF�� 9�ͱ�8.S��¼�2 �+��='f����R�&�A��	�mjiwݗ=/qy��u�0#�yy�o�&`� ��ٲ�|�m!"�@#�g����(6�� ������P)�k��L��+�	fx,x�O3	�B�!r)�ձ/�8��_�!d��.]\c�e����p�t%�d}����;�D�(nv��b-}_���;m}�١.�G<�qm��+V��PtB�49�>��j��t�"N)m�W���VVM�ƪ*�*�D�� �)��
@"�x���W�����n�R�#��/�k_�v�^>�1x
��v�;�˴T|{� ��K�էi7��T��?�Y+���j���[d>=�_���"U�������w�`�m�94i��#Cw�Ɩ���*쑳��t�E�� �I�ImL'U�%|�K�s��>Q�[�|���j}�v�ֶ�]c�'�k����Y�Y���dM�,�|Tʦvas��f�%��h�W������4?�käy'�s����X���7`t��#ॺ� НK��¹Z�yƲG����) �{2� �s#��$����r���v%����ʟ�i;�g���t�IH��H@�bW�̜�D`��Jd����v�eo�E�+�~̅��5y )�_��SvL y�ɉ����O�
�\����;��6�^��~�ן|
�&z{[����leC�Ɯi�I;����
�CP^�RP���9so:�P3W�m��(���(�ړ#�C�n��e1�0ߊR
&J܀��2�1��!�9|Vv�4w'�U���[��ĵ��;��z�mR��u�i�o�ja���xk:V���K_�b�����.��C�zZ�@���,�L���c�{�+c�E�t�꿋��(Q��b�-.�$C���M<߬�_�$3�y�a	��"@x��v<�����>G!2���<ᦒ���^���L��@�<��/9�Z�7�=E�Xzr��< ~��
{�`t2�QVm���Tj ��֎�F�J�.=b�p8��b��P>�g)r42��f��ծћX����kKs�(1�#�>��UM� �/O�m�)Nw&�UZy�:�?Ewcy����t!+�6�X��|��V�i�k����Ǒ�;f�}���o# ��LWĦ�,g6�"��ʽ.1��H��[E/�^=R��.4�L�v%߷�Ʈ�"@d)��u��qa��OWk��j�Pd0��@���
�׿x��:l��ֈ~Tr-��"�qFJ�E�4{[~=�����i��6���s�CD��i�g�u�?�U�*��5�WK�0�?���n����3��ڇ�'l���㐦K])'�"�����(BͿ�p_�o(<3��D��q�,M���<(�N�v�)􆱾��"���"D��?rfY�J'"������@���il�����l�e᝼{����fŃ�|ѳ��JJn���\�bXw���C.���؈<�\���5'��{d�S�R�"�ՊR?�Az@<(�}�}�; ��J��x�$%�y���Ր���Z�-i�]=��G�����B:1��_��)�O�7u|�����ʃ�(��Z7BĜ`Q�jW#����@1[(\��%�ȱSP����;�xO�MWC��vh�~��q�X"~�9��=/�W/��;h���ߥ���<��<e��F��@/�پ�jyQɦ����.�2�j��B��V3+Ҏ�Hq{���g��BY�ׯjϹ9��T��
t:���u���.��ߊ�8>Kc���X�oT���Ŕ���2�ަy�m:3N���"�#^��C
��l@c?X�$D�V�o��B3�X� �#/�d���Tc��o�}}#u��i}�4�_��i����L���{�wb!}��;ȈE�u�̀md�ػ�{s�j�B�MwY�ܖ�1��14Iog�8�#�\t�|�ߴp��$�|�SN�(8]�D2=��"���@�kE�k��岘-��6��j'$�
䰗ZfߦUa�~�����4iXy�R�xs����IUb�Y��94��+���s>��+5U����f�wYdt���:����A��󩔘��sfZ�����/�4��`�(�����k�o0�����t�e,�S��	h�F�%��6�ž��|:R3�<�d���֎�w+��Qv���
MNV���a��7.��*�Xh��LZz�|��H�-�� ����,64�Q�Ĵ���
`"IC���a�&��:�=�q����K���)g�w�|U�3~��݌2���J�)���0w$s�**:��a��9�;s��N�e#�N�{5���]��=0%8�%Z9�m��r}�0��٨}�V�N��,K�C<�s�c���/��paps��ұ3��-؛MfVAV����n�Ӯ��[_�ۓ)|吲���v\��e�M����!c@������)C��\�M(�d���J��3��p�%:�1X�Τ2DN��F�v��J�ؑ�nY�_�Z���AD�r��*��C��u2>>aLIB6�=����N��5���)=|^��Hn�HP��>�<0�B5�c�3��N�5��Q�q*a��0���#G�Qj��l����9�x-i[,_]��uT�r�.�Ǜ��0]6J��<�<QoaT_�r����"����e�:]%.`�d�dUW��"�ߦ].��β��`��T�2� vq���:@�t$^Xh-�|����y�;��l�.��|A�����ڴ��&s�a����U�,l�%��?�P�D����E�#�yt�y�d���Az�=�]1<N�<�Jݤ�ڝU
�L',�x�Y_��l�XHj	���3Oy� ���hm���;�w��2�h�<���kħu��S��A��Q�5�m6� �o�9p���f!��I���U�T�΅0]2͢2"o3N�S5Tl��qa��,�M��$��$�bt��b%<�Q2Cש�Ex�q�l��o�8BU��]�3Od����h�ץ=��B;s�T���Gj�$�}Z��S;U8
Vs�݈'�ta��#�r��I�aWoJ}�/4�g��U�g�99O^��3g�>�]���;ۿ��2�E�t�聽A[�U&��T����~B9g �I,�_�݉�����p��J��n���o�T�O�'����%�{.m��h[̠(� �{J�r>MfyY�j�N�रw���1�����Q��n��"��L�>�W}kw�&Z?V���^��_c���y�W����xV��U�R��:-��7�Ś���r^�^�7���m��S[��2\K,�����c+7�u����O���)�T�����/i�d�y�c�R#O�\;dKA\8M�?��J�Ȫ�3����D7 �hB�l$�����V�����g)^�2*�JsJ�Ir���bq�sW��:�U�Z����_�����0�f��v�s�}	�>ˎ��Y__�D͝#�K��P��*�����$���W|G�/3p�L�۸���YP��-V �d��:��I}�1O�C��u��ݕax��p���hd3!d*�z�GU4>�L&�P�%����#�5
�d�_��8�c1����)3䵋���n�����F�5�qk�ݕ��0���{��^�[�w���-��L�� ���C�C��\K��>�ŮCv�G�p�$�-f,���m	����f��a��S^�,T�[�v����#>�l^�<���cd��[`�	��C�R@yȯk>��{�v傝�3�$z�z�v��Բ4ݵ�B�W���*��8�IY�Kp���g�j���f�v�
�K�/b�-7���
�`��O�Vʨ4��yH/Z��/�^�t}���!�U,<����u�b,��cKz2ͳ�x�/�ٵl�M_Y	N������ЉTbT���M�o�Mp��5�l��m�i��"�Q�m
��\ae�{_ۣ-PQ
�r���'	u�%��j�p�X�g���E"�f��ׅ�>j�覥�gu�.�>Ņ&�m���(�ӺK�#����UǛ�	��J��ܓ��Zk��$��Z'�UQ���xU�_5l6�Ŏ��[���Yе�����6w�>��z�{�c��X�A�Mky6�w-Wӟc�d֙ ��D�~�����~^�h$�[��|u�{O�W���[�έ��+�=�y":��w1����&W�ǿ�#��Bk>���3��b.�b��uǦ������;;讜��ֹ(�Zk�5��`��gow���������F��y(�T�]� ���Jc��? }��/*��6~ܓ�D�O��W }Lq4Kk���4�ae�j7 GL�)B{��ٌU�����,�v���'қPO��]<Tw�����S.��睖y=_�J��]A~��������+B�13?"��Y�fj�ۼ��i��ȔkH�4O퉕
����Y�I&����HE����*5<]�S�����oOa5�u��9�e�(�i3C|��2�B%Y����gWm!'�>�MAgm!<\5tS��F*�A���Pb5X<>s=��<�9i!��B<|�c�/�g\k�[t#Z�n$��f�J�\��hz���M��>�TއڤX��cY�9Vܟ���4�Ij�b������K����_ˀ�B0�e"z��� ��`4���.�6���x�l�-�s6y(��X�����Î�� �_��x�<�M&tXdY�[dK��4e��C��z���(��
{!�)����P��M���1��*�:&�]�֜GX��S0�ңj�@��3R,M6{�����S,�+{.`�RCيk�)O $D��%zp�kfM�a}BǨ�nI�&^&�W��N��-�M���H3P��)n�kr0��PN�>�z*%�󒿹t�A����錦�S��������D�z�i���	E����ѳ��eJn�G�r�]m㾊��5�GZUgBC+E��N����>��ڈ������ձ�_��P�DN�p�$�pOb�.��g�;+��nr{�G��g��4?V9�pf�lGݛD�R� E��_@�q��"�p:�gNkI�:�|O����a�W
�I��$1+"�r{sUú����T 80�砅���;��H"��YC�S�iYԙ�PeE>�����P�5��)�k`� i(��G)���ҏj�E�L�o���fϷ�E狋մ}wI�����J}����!4s�������1��V����(��i���w E�l�S6��Ԍ�f��֒�Ձ�TV���+��}r���!�Et��Vs�����9$���wM�@�&�4��v{�Y!cI.3��ܵ.�s�F���x1 ���J��Ƀ��I8G�|��ⷦ�k���Z�%��_�iO9��p7�p�D����3ek�;�@}��Tn�!�\�a�&���ʃg-�	��;B�J�� 2f�-����Bd�Un�s:�+�<-���������Hd�KPܿ13"�ܕ�r��8�ZJ�on,�<��`8�r��,U��%%YK��#�- �suV��N��o��X�+Y(J�,<T1��YX/yR!^�[�v�NPA�{^4(���=K�9���ԢZ��h�Te�TW�-�+,��h�������j�b��Q����-�1���k�.AF%���i���$��/[�gǺe��xݺ��E��{ɓ�.j �D�f`X�q9�����e�en0�ʩ)Bi��P���c�H(���J+�����֌T��N����Ir���~���K��{㳹����������GT�0!�ɩ)tq	vZ�d��xO�eeˣ�t�����T�o��%R�Շ�+G���8�*�bDV���b�%����zR������ ����K8�n��Rs.*���v�4�Dt��"���ZS���]^x����{��hj�����1�Je:{Xc��/��'A�ZӉZ��w���B]��!��L�n��B#���'��N�O�VZX=�W��b�A���;�pB>�6 ��~�q�C�#n� �A�N
�T�׉mY����(?׿���J�Eob������̗�h�%B��I�K\��	�^� ~�&N� � eF-H�6��k��8����aR���/\��r���r2���I�E�����ߩ`2,��.�1�Ǫ�.�3�g3��=������ܱ$�C'9���PU�#i�i0l2�֧v!�!����\m�?h���;L���c3��=Dc����`��h���WM�P�sOQ�:]���H��G�5% [fS�9_zC����h��5�s�0��?�થ����ބ�i�o�Q{�>ʁ�\@�&p�ss�G~��o�v����O0��u#�� Z�T��s3:2ks��K�~�����x(��v]:�q)��Ⱥ@ߧT:����@��h͏�ͳ/+Ym2fo<�г��3-�*���QT��ɟ�]�����V��V9�J�f.s�ZF�6���,� 4��j�t�*���$j�+�P<�J}"��3ÃZ�����rs���;B�%dS��>Ϗ8�ۏb��f��ڀhu�3R����S�ج.��4V�R�&o��MM��l>�;M�����櫤�-��&��ƴr�cv��S���R�W����*#�jG+o`� v!P7V�7T�g���V0-����7&A�t�|{�},��9������ nDM��n���:r�E��9i2X� ��ɸc�_(Gu,~B�$(����xK
����y��{��;?:����I�k��NvAt����\��y��$�G�EX�?����H���'�LC����
Ac� �m���$�"�Q��0�e0���u[O¾9�Q�z����F��Vf���F��A������wh_��Z�Ў4�ʄ��,��i���'�} ����v�r6�M"������gj�9&��5�y�>Z����:�î
`��r��)���)x�D<7���qgZ�1T�H��؃��ф����Q���g2��y��u�Y*k�+�ǟ���`�/$я�����d���<B �6��f'�Lʘ�]m��N�9b��e
��O$~�X*�-������a��B�!�
L/&2Xf�-��}���R5�� �)`H6�,2��x�I��k���w�[3�ZCJ�H�aG6;B�e%����)Z�L9\B{�tOIZ��:M�9�2��D<���Rn�(qX�_�����S�%_��D���h�����}��켮
�@p�@yO;ɮ�NJ��߶-����̧D䰬C����8�E�i��JH0w]����*{$Q=r���3X�*����8���p�l�Z��!�3]S� u��Ck9�qZ|�7��	Һ���ٔ���67��e���Ɖ�s�l+
4�+�]�h��|�^xkW��xr8B-[��=V�c�~�^7&ח�P�6ɍ��Hhu�J#]7��z��)���}�e���&�&Q_�NQ�&xg���2e�&g%�ؚ/^���v�9��T�<O������곫'b'X�V��n6���)j���j�ZN�*ZOP��^�C�~�~����2����H"�ay:�yv����� ��C�t?n�"e54B}g��������\F�b��;[�����g�b ��w���P�N��vT��m�~�(p��+*8J�()/�I��=�\GQ븈	�̋l�,-Z��%�M�fT��dEv��"�_�7+Tj�(��D6��́:T���B�Fs迮:�솷��%�5]E��E���2>I �>� TM�:�ya ln�qX7u �jOu?���-��K��(]R�ܽ�y����T,O�|�r{�h�f)���o��ۂ D߀თ����Y_8�aٞ��#+��9'}��*"��*�j\	Q�u�+F]����]�%��U>�7���+{" �B��񰰠���.��.C�d��sM+�L�} ls�-.q�d@�߬(�i��������e%�X,`���'$Q�����(,`�~����Uy�e"���P���4�?2�`t|�3������k)�a�� &Ԡ*�=���F�5�tq�:Ä�_$bӘ����:��W}�Wr�gE����\6#ǚ�|�;%���j-@�Q�1�맲7-A��NAs5�4�!\]��s��l��Vx,&s8ptĄ�}�͵�EƔ�M�ڀ��vD���3�C[��W�C�:�Z ���|�����X��'x#m�;���*�u<cGc�����1�bnh4g�PHl����؃'�Ll�^��sԛ���������߇�lz�8���uU��Άġ�����wJ�|�פ�'������j���Jj��N�kM�݌7ǉ�S�����m-rF�W�(S@�W?��ŋ�L2ԯٙi�䂗	������gD��v[�`�x!��Q4�*�^���w��N�%nY"b\���a�a���s�S����q����[m'n_`���o�i,͞Қ��}�9�^���ѐ����+K8u�
)1�<y�'F[i��|���#����̶oU��)>��"	鏜hh��j��\<c�I��4/�r����^�8@3�!g^���餚�>ZH��p�6�l�	(4U{�~;���HG"���x{̞6�|� _?x������T�p�D�X�5�Π�|2��h�%H1��~����d�v�x#^��g�1���Z7���-x�bw�y�D��]�Ǩo.�2_��(?j!6k����z�q�*W���̨ӻp�s�����QN+���Qw�|��á�"�/��[���z�7�����u�K�9vm��J�K��Òr��۝HI�P'ӝN�-��U �}���Q���N%;��C;���O#�ؒ�`��*;���;M�&�'�A�Fl��	�_��d�����e}	d��⻃ą���gjeU��*��6f�E	����T���i��lg�R����튚C�h����6���+z��n�Bz���~&"Rf�X�$Rytʡ S�?6b-pĉ_�J���}�Z8��fOY�Q�r��lΨ���5��T�v��8|�"�*�������SA��8^d�))G�<S:�%^����7�}P��J6�-���;������J�Qe���1b��y�/r8���|M�7#;�9#"� T��0�� �٢K�r	%�9�y�h�~���Z�O����<�K���\����XV5��#������g�W�JsE�f3����X%���Zr��-����O]C�A` Z�A��!���&��iR��x�B/�E�ҝ� #X���>����?vV8�,F�^e^P[v�ᯒ�oOLLλʒ�T�s@�L�<�4�0�p��I��dQ�}��aUe[T�v�7�]>V�1�,�9�!?�2�����<<D�$m���:s���OQ����K�O�'�n�t9�`�AJ�m#�L�l�?��3��A��po;�Ar}:[G�3��o@��N��="<��=s�� ����/�<O��NQ��)��1�z���.�8��:�Av1%&���ɝ�g�:�D�ށz��׳^R�������\C�#,̳'縇��Q2�(�k\����jPLO��`�����øK�Uyx� m%�(��@:4���|T�.�|��2�P�I����)�)��]�� �O}��|�1�ʚ��"���'�kB�)0����>;��!!���s���S�HP�QR�]���鹤���hʝ�kb��[�u�F�'����6 ��Lt�0��D�~�U���ω�����ݼ��w������[	魃����(o��[��ώ-�\?>�P��Z׾���e{T7}e��K�l���H�+K��S?�=|��Lt�v\R��I�灯�i�8�妼~��`�t+N ��5� [�����-��wl�G�� ��5!#��t׉�U[���Ԫ����Q%E5���鼔	b�0��1n&I�����n�=\F'��]d�+.�������\<���~J�yV�H�)�%��6������;�o�M޲V�&;�.%�
	����1�L`8�4�
t�*�w�Z/v�5aV;(���`, x��>bfZi��#�s!���Z��8��f,9��{*�q�H��~Ex"ѴT��c����ד���D65H�I�Q�w���C�!u�]���zE�=}!ɨ-��1�%�i
��@��IM�t����x�	����ޓY�\����"�j���S�ĥh۞�����>�12>}R��)ܑ�� ��Z��t�yve��'�������lٜ	zB,��N��x= NL�����6c`�w2j�>���wE^�U�����mcz�ݵ�J�s��'�cN9du�-��3���E'�#2U�P�%+���i��6� ��M���֞d"c���Ŏ�AЊX���[�a�lG���߻�G ^ �Dcsr-���R\O�	�i�@��=e6�9�w��� ��A��4�a{ؖ�ݖ�|o9�Jk�z
e�ѽj�xY@�wR1�tMa�6�X�}oT�SV��q�R��[.�k��ͥ�>�H���m,k����� u�6�z�Wӂ��a��4m����Z�:]��Ѣ[/]� �T��\�&=1�	k�1�:��u(=,	Մ��(,��cN�v�\�����"C����Ű�~9�ԝ �{�3UW�!�i�p���*�c�9y�S� :��}_���`t�G���i?��۟�P���f��I ��kw7��P��9���T������Zd�j��x����`�������2�e\�bl�^�����6���<Y�l5�l�}<��);쒊�!3-��JW���|�Mi;R���u��싩7���	�M���'����>�ې���:O��V{%XwhRh�7��W����hj	�Q��1"(�[d]�D�!�l"1��t����e��O�1��)O\��9��ܪ@A=��m��vO���pR��ܜ+��?ͮ���R���6X~ҧ(pQ����L�@��tķ����7�=�u���QuQ�O�o[�?�o��H��ϱ9��HY���[�� ����M�`�}�{�I�SjD��!g����Դ��K�w	W�	d���5�C��.ma�!�wʢ�y��{����"�͐�O7U_�ݥol�����5��L�V����u����4�-�̅�|u���q�r�V��AW���DBҗ(jv���e�c�Y,ۯp?G��{n�� ������-͊�v���!�Љ@>���%ui� ���=W�oǲ�eK��|�7��)FR(���?P+o4\ Z�Pc�A���|�J0-�k����N��߶���UFH��;��z��}���~S��M�����S�9�$�$�� Fz.T�* 199�� C\��f�b~UZVW��Ss���|5 �Su H �f�H�[B�@��ޚ�.�����F���W�Hv/�ѕB�
ZP����^ŀ�&B>�wPM�ޱI�wr�Ԑ���v�88Ig�9�_Rm�I�[9��+��*�BHoW�U��ɸ�t$i�!+� ����e�I���v���C�iK'�u,*���Tr{cC{�����"b���`0^]�u�^^_��n�NMT�Ϛ�P�pƝ���I���|AFE�W��sJ��{M�;�$�o9R�aR���0|��ד����{&r���_�E�+7��Ŋ�{12/������t�O*"�5��eOZ�-p��@��)q����Ҁ�\.a��t������IΤ+��L�A�ȑ�*�|KEY�{D5�;rI�1��V�ڏ���[� �0�]��z�9�ڔ�>>XxsF���J�����L0F�/����k5�^ �e�\S�����~�m=s���U��;FٔS�@L����P;�XOY �.�y�Z�~Yv�˻{��$,�l8~�@kv� ��A�������'�!�6�J�;�L�$��0�{Uh �EK�o�e��jق�o$#�����݈�}�$�/k������\�ђ�	h��� P�Pp��\��,F��{ ['�CW�oOSyCb�e.)C�ېh�,�Z�T�?`������}=��X\!��5��h����uy��Kuz}{[>��"�P�S�a������	)�>_�S ��G�R��x�gd�;��v*A�@V[I����̈́D���Y��&�R�i�W��������t���v]-V=<V2��:+�|�;.��E'��ѵ����Ѓ�BzY'�IY ��D�7r����OO�	��l��
t����C�YX�Oo��@�J��b?m�� ��|0�!��\�{s���K!�pG������}6�jJ�#�!7�!3#���Uκ�:!@CX��^xO��A��;�}X�> ��$��dʙ(K���7�)<SG籆[�D��2� ߄���k��X.>����שp�g�eXD�V���5���ʉi~H��9�
���߰ad��j��|��1{�RcY4S)��d
��Ƕ��{ef:]}�W��}�J�#'N2G�0�ٮ�|���¡����g�8��mK{���8��9��*U����x�Jp�`���G���h�Ǚ:�Z�s�D��y��P�7���vD�ɚ�*"2���U]�4�E�u,^�Q�H��)�M���|_'�Mp�3op��AIs%�ă(��d�����w+xb' �I�o��6�2��D�9^�T� �C/��m��qP�F+��� �T�`�<��F�d���;ۯU|�5�ZymU*X�`@����{Uώ�/d �
' �5���G��م�'�4�U5�0_����o����Æ�
�C�]�b�г\����|�1���N�;�#l��0�p�X�{�n�C����>�PDA��8ܭ�|�c�_@a�RO��l�b��x�>���
0���,��n����vT�4����.v}d�G���2cm��Y��)��ّ�7�g�� �m�p�ÓR���q�_
�aԖ��b�c�'!pe��Cًo����
���d����D,���=n��GwF�Dj;֪��T��P��gp��@�?�D�y�'.�:�Qu`p�S�ö�hC	0�eA#�K��%�7t9�R��!�jWu[��L�?�/���^��R��൑�xn�p�����L�5O>���uC~WGZI<0>PY�W������#dpG߯�J����e/U�7�/l���7��D�8��V#[�ܙ����ɑ#���坅S�f��%�ȡz�����$��b��M��1�d��1_M\RG����q1�(?�%�T��Ý"�q����0���i�V$K���ϥGg���O�}9;NIi��r%�"Q��=@*^�w
Xȋ�o ��<����ϲ������=/�>L���}� ]	*�jU���ֺz�o)�NCt���=>��,��4D�v`D<C���óe�+i�
���a����N�1�PN5[����(g%�'4��i6dDV��w֌짢�e]R��%
��g'�F���ߢ�k�Kv1��O�j�5K��>�*���M�J?n�����2na�;�%&0뎡��Rh
\��M����B)�J�o�+�_|�	��Is���@`q\��N�S;C����uj�]*D/�n��Z�>��j����$�)+Z	e��37���I$]>��]�%�4JsT�2��"��\������h{N���X�]�"�]/?�Ꝗ���0�1�Q�KO��6h;c��3��6�a��A���eZz� �8y\��w^�}?{͏�׌�1�9����A��ȉo8Z�׏�Iن�vA��vB�� ���X�_[�sq&C���tf��2H�[&��O�[��W���E�#��s�/#��_�G��2f�4�z=�+�{�����D���y���������8tk8���j�Rm��+��m �I�b+ԗ�}�)�mͩ,"cy�̀��_!�Ҳ��F�<�ޜP�Ć@�;���BEױ�0Nr�dj�Z���ؓ=���$��$�i<V����JR���ήs�ކL0j�Z���ZY��~����#� 1e- ?s]�7�����~�=�[LJ�mc*�O��<� ��Ї��<_��.ˌ4#���-H����b����a���ɬ1(֓X���Tx`l��9x�U�]�lr��	��ۓ}0�9��N�bӔ�����n���7�3�~*��4vM��~�z|uHZ��_<��y�z���*�$n��S�?�Q��?�zy�x\�k�vϓBǏ�!�\�3������ZV��.�0��Zl��L�E���i˺W���ܢ���K�,��ҋ�Gs-/��@HB�y���rS�aluZoңA�7x�WݯV�xQ7��,a1\�.k@	F���;Y��lѢ�s{���^��@2g54���M!!�n�b[쪯u��.g>���R��9�p*��4X �& �UӚ��{��,�m����D;.a���r0���m@Ԭ�9h��^��҂�D�@��5�*9�@[b�Z�_pШ�O�`1Bj�	��SG]���#;[�\(�e�5�9�����H;o��r��v�b��N�9��{tq�Ŋ�eQU��l?�\��Lk%����c&wJ��gH�Q����j������ fE�Wj�ө��.UQhS{��^�E21���kK�����2��7�����4[/<�$¢s�J��������7�Ʀ�6�ٝ�=�+Ԟ���D���X;��l_[���$��������Z�X�b�Ld͒r���Z",�<�f��a&gpg���v�R�%��cB��t��&�K�mz��� ޴��f���<f��y�zW�F:K�~���"�-���;�Tҋ"Ȯ��o)#��&�3���
2n����0?���\���B��j�ƴ���a5��	a�yL3��'9;ݴZ���<lV!�G*ߖ�G����V�r�Oīkf�2p�tH����]�rh�ޗ�v,6y�Ǔ)A�L۳���|[�� b�(�.�j����;�)a�5�a,��p���� <�wa��P� ���[��E-���5@��޲��M��T���x�o�9���]'�2����G���Ձ��Wh����2&8���[c�2����(k2�>��0�d��,��/��2����lN�;_ɱcɛ�H�ߋI�ˤ^U%�h��	L��* l��?�2���QW�m���]�kx�ʤ \�<�]W�\55�+��]~:\fd��+DX�����{�3Z��f����h��y�%��w?��[k��D@G󓃞x����lU���|o���#hZ�H����t�c4qC��A�H\$��C*`��Vb,���L�m���¦4�.���+#ҝ��0�Z�o�$0r���&fb6�K�8sR�(�[L�ҏ>��n[	j���9�&�SN�!1����MC3�Ftc诰r�i���D�Q�8w�N�l�I3�hq�����^��4��Y�K�z��֭	 �1�
���]�P T�;����]g'_��KS�6yTs4co�'���1`���6�=j��AB��=� (E4��G	4~� ���N�DhW��&�h�/E�U��T�qR����졆c1(b���翢XrK�#�x���4'���Ψ%� BK�aX�$���P�W)����4����෼��.l�]��#{�|XJc6s@�9�nk$M�r�`��S���7:6���z	���H�!U�(����e0�8t�jE6;�!��ģ��.0;���A�P:��6B�Q��*GR��!~��(A�Ա7���A��̷�O�,�^C�|�p���R>�,���(j�*�~��`y�UU/�Jغ$�ĹY�s޲5i��� 㽖Tl:L����D�֎�#�ͬd�$i��i6��5x"[�q���ׂ�:A7ĮB�+�Ǭf����/{�F��P�f��������i$4q�V�u9�&�V���h�m�M|���p�kD�@M��	i ��?�$�A�	����O5�εR����d%��ȏ�֤�
��`������qHF��EK_�I���5�c�F]��R��P��O����5_�_�!3^�iE�Gs!8�R]���ܼ�NkY��jij'�	$�H�����D�A�S*w0f�0)�L��Ow�[a����9�#|Es��B��'v�{�]@���0�p��q���ȯ��Q<M��N�M�3���Ӄr�F�����y����A������a��6�\�=���#��,A��:$N7�v/�n���*����y?�)�4$&�θFp^�kz�鷄k-`��y���H�fnI� �b�"�2Z���\���D�U��O$~?\��_�ft�FV!I��m����̇
Y��s��Z�Tο,����HQp�1FKg�?]�p`=ݭȢH�n�B�Z}�Z�,@U����gg��������.R��*V.*��v�n�wV�/ #�ץ�tM���~JLI^Nb���z��ly��2>J�ҍ�{�u���	V���r�Zl`���4WI�ϴ]++�VJ�� /�9Y*���Ur92�56�εX��Љ��o���Awt�_8�D�ҁ ���a�g�vI��['C��Y�3����~	�;n�%�S�U݇�i{�����팕-TQ C��d��������%���1�W���:������3O}�W(���U{PWXơ��(�c�G�j���G��ϭ��B��n�TO�����ޠ&�A�NS�,8	�y:=���������˔��{�x�6\L<E�x��z�*Z�qj���"��ت7��5ktB�Y@��kL�g���8�ʊ�������J(���	bߥ��s�U�ՒBA����k�["�
��m��뜎G��5KNͪ�2�-�_�g��_� ����P+Ⱥ��C*�{ٴ�F-��)S�T*�p|�X����BD?t�X�L2{h�p�?���kM�i"��ĝ��g5�1�N~8n�&z��ï0�U��`꺓`�K�D�lZ��2�є�~��c�0�OEf���w�p��: Qrʹg���S<��W��xTeH��9���f
���\(�?�i�VB$8��{-�-�@+y�S}B����Cq�������7����71��}�Z���k]���ѭ������K�j�sl�y���%��p�q�c���	r�u}F:�iR7ƽi�ꇳ�1��j�?�e����.��iӡ7���}�$�Y>uD.���$_��%V���W��^�ܐ�+	P`�W��]]?R:�3]q_,��mh���}�N�d~�w�~�Zt?o�k�ݳ[4w\���@Ty
��+�A:^�臇��2���/C�|����		�:�}��|��x�D�B
Сs��6�r1����)�<X�m�,m�XKCJCR5ro�6G���jJ��cDo�Z�v�H�}pݾ=-���*k��v"hW�������~���5WG�<u��G�Q��vۊtQ�>�7�08��UP4�-Hx^I�^���-��\ԲS�q͋I���a��,��:�~_�aA�����jMéҵ��L(�c�E���]��g
�ެ�0�����L).Oo �"���Ȳ"���QHҐ�/��)Ц�y�+�{��u�����N9��~�����te�L��[~=U)�(͌Q��i�,.{�`��;��������������!��^o[b���+Eזom��L憧f](�"�Q��M
Km�@�d�# "��������{̡u�+d�{��/�D{��j�81"���C��ν����m��,^j"*�� ������p�U@o��!��/z��N<0}U�1�\IV'�ζ?�u}MR�C���Aw5�*Y�����k{"�ˉ��a����JO&jrvdr�[U��N��
k��.����D �na-���s�3��<F��}�
A�(�@��'���9�_i6+����u��A! {0r���&�%m&��܀��I.g�_�F�6���T��(������������^_�݁���.��>���ƒ�Q���o5��w4@5��-�q�5�i0X � ��oS@�B��ח")�o�Ev�/��Ѐ�ŜE��]�7.ͷ�� tc�gtD�ge��9�E1�3Ԁj�M�Q�4��c7�A�쾲d&.�Ը��ǝ7ҏi�L�*��$)�%����k�[P���t�G���N5q�
@������f �q������B�&��b��M ?��].�@:i�̨�Ѯ{7�����T�[χK�-(��>�|t��r��ꒂ�䚒�[��c�6	�H�	l�P��K[����ty�6�gg�� 3�!�8X���'A=�Y������T������+��
g��7^J���I�i��OQ>y�?cro�:�Z��e��w��ӮD�],&b �>Hha]g鈫䖰��Uұb$���Qn^�GT�������tSُ5�d��[�X��НE�"#(u��%qb�H�GJo=�����K��;���e�N��x9��|S��*�Z*Th�0��i���g0��miG���IF�W�/b5(�	�����
����;'��2O����C,�l�Ѯ�0�U��M�t��7�а
|��{���2>�,����H&{�	�%�WT{�v����/W��L+������|�qȆZn�l��^��b�ah����p�� �ع��n�?��G��uE�^ڼ��w  'U�g�#���&
B`��$��.>x�m�@����fR<x�4����c>9�n���PH�ߎY�"m+SB�My\fa�������,��/�K��C�jv[z�O�U}o�l���1j�yBDm���4�W1�#O����5jݸ�?�͞�Zy斸XW檁Ќ}`�G�����t�e�$�3�ϕߌq��?�r��A��a�z���/�H�_�lk��� �G ��s�xuݖ	x�����t͸�هY��(��<�7����?0)^�Sz(6�$j�t?���ry�V��=�C����D�MAj�p�prs�(�Q��F����ɹ�(�y~Y?'L�w�$�u�(t�{�T�6jK��E��7S�v�D���)��raPT��vc��FFQ��մ�F�u���D4�!��!��so-&>���7���������i�놩#GD_�rT��j��i%[�97�J(Z�����S�+�PH���cp,�\��R��a�'ݷ�t��|M�aB�rW�6Q*�@2��V:��ѽ��%hL��z6�Œn��"@;"���T=��j> �_������g�X��;P3*�<�W���&��3��Ω;���l[� ��SE���?3=m2�~�˅UYs/ڥ+61R�%o��ߓ���{#
�h\c۰>�����f-T\&�nK7���ab�p�*T�����
��رZ{�}��
Q�Y�H҉������c���/W�U�f��_?S���硭0��~q� #5��jk�6���ݸ.�h�A��9��T��5C(Y%��,]�$�H�q]�yoi��;�0��sl�h��D���T�$���;�4���yO:�(��1��NV�\��<��t�͹��tB�{�~��=ӝVz"i�<-����0���y���a��`�z����;c����Ӯ�AC�x�l���>�^��3��|;sv���mCJ�Z}�ω������UW=������:��_�֟�:�.��ل��w��i:�k�Gfa�n/Z�..R�e{��h��ڿp��h$0�3/p����*�K䑁~�/+le!��:���)Q!Na2.T����]���B@�\ݹ;�WQ��"S(o�/${ޛ�L�����'�jRST�I���N-xW1� �J��8���n�&��dU6��S�ѧ�fjɟ�+�@���A�9��;	�u-�d=�]��f�Q��ϕ��{���!������I��������nAb�1e:� ��,H%9<���f��<~/-�߶�&<�&SN����8aғC�8��I&�&u��\��즼��4[�*�9N��
�sz��&����]vC;c]u{f"���Z���ά%k7v��!]���!]��Zs���k��mj�w�B�@�tG?d�h̋^a6��Q�ٶq�7iZ1㐵�%�B�L�1��x��ïPX���X���6����?��_ST����ܭv���M�j��C�o\q����s��J�����Di�n뼠0Ĥ���%c��S�3��@�N x�hY�M�����#%���K'a�g#�זsf�q$UU>�ڬ�}��KO �5�<6 �df�}An�^!ŵz	<7Rg�;>dKm���rؖ*�c�06ɍ�T����#|6\x�%\��Ql�Kna�-�ћ)&�1���j�4dM;�2�8�������b.��T�����з�@1t����F�۹䠍�<��e�G#EQ�1Dz.->Z�N�����ǔ�6-��'+J&5x�!+X��z`�(�"�a0�o.�w�%$#&�n�X۾��ێ���ga��cHH=��58ʟ���ASޮ��gr�^G^%�x����.�J[Z�j��.4]î&���+|���ڔ|��,�Y")�����x�x��9�Ϯ'2B�e�u+�� ��2�ui�H�������\.���$|�������m���k�G�j�!��{���҄�A�,r���H�"b��Nn`^ٌ��xٚ�DP=���AǨjҫ^�}�H�"�"zo�rm�a��w+c���-���2���۵�[h�Z��#.��M�k4�J�xA�᳖��,DÀ��麎�}9S��Gئ��cs�!ы�	�O����8r,�	.�"O�U�����nf���8�s�]��q���<J[��ݠ�)�Ųec2�- @r���x)Ki��m�����)���BԠ��z�����n�d����fT���@�\lu��}�-#�`�s��$�7��[����g�\����p6�-�<��u�GиT��>���D��%��R ��t8w{����"�h�3-�o�ċ+�:���h1��B�^?�z!���qA����ܤ�XM��ͮSA��3� ���j�6�9�7����,�[_jB�Q���ΘB,E֕�}�醣dR�\��1ƛ!��zq���Y����@[�FI�6&�.�K\��%VV_r��w�j͚���Y�a�!AA�d$�Σ��9P,=;�;Uo�!��������(z����&�#���|�V�lJ�;�����L���r�*x7�>/	7N�:E>�Yw�w�[����ŋ�9��zQ�Lݒ?�W�cy����9���Fۯ+����%;S��2�uV�V�>}�D���^H��'<���+?�갑>
pe���S%NE4���ɩb5cDȖ��|"u�S��>0B��N(rJ��x�"�]Q�B���Q�b�'��矌�k��5h3ky���U�m�_ �_dN�03��$%t�
HK2�cO9�O������,7K�%T�L|�^�V`��<��7;�E��t�W������^�tv�vz�#��?�95N�|Cn�U�tL�ӭ�4s�ޏgH��ŋO"��#P��r���Va-rrx���I�X@��l��!��l/�`�Д�G{6uX�O�г�ຶ"����/|�I�V��v����}��{���Ҵ'A�����P�������L�l���`\��b3�e�:f�էu�wU�>�;;��`AyG�\�=$���2ȃ��osp[D�/�:N��Y���{�S�q�]�28@"5�ݚ�Q'�֍Q۸���Hb\Bċ�e݆&l��|��]���\V�x��)Mq���c�q�%P�D�!�:��"OU���8��M�L\��i�@�95O�UJ�k�sG;;Λ&o�&qP\m��=7g�uAE	P�dk��7���I4ػ�al��
`�~&�l�؉�=�(y��N�_���1��f�ߛ��Grrr*ōf��I^��v��K|��~Our�kB�Y�<��A4g��;��K����=S^3�� �4���L� [�C5]8��mV�J*��\h���`-gޫN4�b� �����NNDk��͘7p� ��mt��NL�Ĵ;r�㽜��Y�m�P�JEcj��.���Ԭ��1�਴Ty�e�����]����&�u�����ʄ�B�g6�1���W���]������>t�.��7	o�7�	ɉ=z��fv��f!۪��E��)��93�u�0"�b�"�Q8��5��������
�o�;�m4�;�f�4���vP��|��h.4R�l*�&c�Ә4{�$l���w{	񵙳��ަ�
�@�ےZGI�j�:����}�	��N��r/�C�>@�#�G�~r���w�=�i4摑�W�P��57��q@{1�&������!�-�(RWoI������=և����;G���<��H��x�����45�N���`H�A���P�o�����}�|��F���I�%h4p`"?�������n���E2~�-�})��SЩA'���[�	=9Eh�O�]��vn������g�W�P	���[N|�n7��w�f~�!��fy�X�&y��R������M����\#O����QD�x�E�i��U[s�P(¥�����[�F&i�k�
�,3������9��1D�RG�0�'��+�M��6�&X5#腢_u]N�I�Hob��ߡ.������wͷ5����gk������_#��v���B�8#�!n���g�O�mE�YOY����E:�&�-���/� �u�E��IgƠ���+�f�N��N2 ��A3OUTF;�K�܆m�s�^�@���;��Q9L��T/��JEb%�ė� ը&	L{�s�$נ��]��]��Z;�>F��E�dͮ�N$K����ο��[�n�8��T:N���2I�FI�!�>)�vo�����&:g|��_�g{�
��C�?�%F��2���B%��O2�A�M�\���%P��,sI��n�;��u�n�L�Ɵ5�E(�I����ƜM�LϹ��o�1Y��!�&~�w�л�g���zT��5��t"�*�Ex݆��ȁG4�޹�h�݂�(������6:�e��k��}O�S|ݥ�;��K	�@�h���}Ҟm�"�{v=�_fd-կ�x���gȓe��W�)�����ei�C�O'��4�3�����C�H)N	�kZ��	������/ L�^&m�ky�>������/%r$GYR���ؚ��s��� YX]za�s�A>�����|g�� �����YH��js�`�^���^\�=҄mw��B��:�V0Bg\����ׯh�l�li��6�9�`zq�
�W��$m;���FoB+���=�F�J�^6��v�,��3)m���"#6���MlY1ޘ��PMz��	�n�жE���"�{���=�'�/�AC�"��d:��"��%N�4�><)�Viܕ?B��Q�7c����Zy%w�[����T��"� �)5�Uԁ8���<�0VBܑ��ШŐc��{sd�z#�T����bԂ.�� �U�=+ƭ���/L������+���i1V�� ��QOVcgҍ��e���nB,��c��<��K�,A�@��ӣB2Ul���`�4|��i^9il���x���ϔ~����'!Y��n͂x޳��=�o�вNa+ΡU�<GE���1�O��a���8�)��jI��^Oķ�W�������3�U�
�ڴq%��z�m���|�֐Բ��M�m�?�EY6���L�	h��$���c�=ʽʙ�WGx+�`=m��7�#]�R������ש����`¬�R����^�\wa�nm���͠`5픀�LKY;6c�PlP�%�Tc�|h�U8x|y��6�gkשgT"�k��e�����=a0��`���f�@�N��P-Uda�(g25l~����d<��X�ٞ���?n�39�������y�@�T@�ͽd�T�����9�"R�P���|��>��W2����&'4�,� ������ҹ�U^���Nd�
zi���W�� Z�j?��<"�������+�J�GS�4�j����Ӭ��	O
� �{�.��h���F���k�#�X;�n�w�0s�6�,z�lϝ����D��}ũg��I��9��W��NH�3;m�^"�~�FdT�ic������-��~�9�2'���� �QN����������������+>�ƴ߷vѻ����)n^�+�T9]}�bw����{���9|�4�Y61�=����&�v�0?������c��}^�z|�ӽY|Ysw=F�[��'��|`�K�;#��nƾ�1�?�0!M�� �r��{�D�J9��?B(�9S:�6?��O]&�8�Q��Rd�Z>���v��}�{��N2�$X��bƢ�yLT��T hP_��J�e�f���6���/��^� ��Wɐ�=�̰�kY�ĉ�[8��1iH.2.,~�dv_�$��Vc�H��%$3X%a�xs�?���P��ȯ8����f�L�f^����{ڞ��?�ԉ�r 5�&7μ��2�I�HƎ�<�:�m��C�6��͛�BP��D",q��Rux����@�JY�f��
3����%�3Nu)
��R�#�
a�՜>�E���[���UA���҆����n��%��w�������ג��i��Hjr���w^�\rx�8O���s'�� pC���^h򚲟��>���*�0`��CZoM�6���zCr�ل0Xq�
����ttiaݰ�X�	-��U�?�f�i� @X��>�`u�Jǥj����zO±T�l�9AEиi�C��Y[1�~$+�ļ�@6.�棰���N���%E���L�}_�J�6a���߫,�}2�0�i�܅L4�F�:G�l�LT|��/��g?a�):��A���@�`���3p}<,zw%ٕ�K��[K#��NX�-��O�O�@X�m�mS����X��A=�.Ӄ}8����n��M��g�#~���,>٨��"V�Y����Hɉo�y��!�q�|q����j�Z����3TU�2�vv��p���m2@⠹=�(%
3<��݄�pE������m�ݲ]�f��J0o<�륅(H(A���L� 1���.(כ���i8A"����U�#�l@�QQ7�}%ZD�{��p��т�{�,�ށa��Z�'y��J#|��WH0t-�5��$t��V� Ý��s�U�FW��&�!��~|��E���;1U@y�qY��oZᥖ���@�t~��E�+T��`'��1Y��]	C��[���S�5��$�2�`�6h0r��3�lr���/���9rJ�r'{�Z���}��PS�Xu��Z2>���ڀ�.��xR=MJ&Bg�դ���}���(ә�,�V�/Y�"����J��5����4���v�wͨw�Z��0T���C�e\�c���vM�^.e�����Jbc�m�̪��fۚfW;�t�N!a[���{A�4MZ�2I�\�|�u�X	%���GK�u�^��=�1o�1kY?T֝g�P'�'�T�p*-!J�A�]?R�X���x`):޺t��e�̺�&R��� ���7p&\ �k��"\�{�'W= +L	������ˀ��+_��;��'��E2W�C��g[0��=R4���)q�N*���<�Vp��� r)���O�\�X7�D��y�]�u|��A�hD��?[*ՠVH�-�8��� >VL�)P��4{k���Ń��b��/��;�#J������ܙ�:�g&���HS����/���T�U��#�3����L�������v��}þ��V�~jƊv�����͍�E�3̀��k)��Q��I9�|1F)`��@"4���2����>��?��	�r��b���7rKJ?�Ẕ�A��|���o�aJ��)�:a�pޛ-�}�A5��h�
��d9b���Y��p����l�l+�B�vK��!Kd:��ۅsxtJ0��1x��9����Q`��0�"?��pB�b5�E�a���k����Zʐ�y 1�H��v�IO�������-/��4%��J(J���BYH5�i�����^d���u��d�p���Z���x�׈`g��`#��MΕwa77���g h�/�<��Q?^	)��Ƅ^ײ��p&[n�����HhA�8ي�ضs�h�����'	(��McڝKD��+҆�7�0�I�7�ty\N��}�\���~��4�.��izJ
=?��]p��JH�j'R`���� �h�Pϻ�qB>���fs4(j�3�RI�a�id�F��˹���Yd;8!��}���fj����KjY����ʵ�W����|Wu���y��3a��Gͱ���I�������P�����tS=����V���	�pt��H7�QCF&�lYg2���c�]�����U�7nհ�Κ�d��I0�(�_Y���k��Y��v4U'������c<���M� ���@�q�Z�'*˩f5w۾s��Ϣ��i��~�c�ܢI�*����o������ȕ�"���z����ͬ �^�������֠h�b1י���)ͺb<���I�$'@����E�*�*�����A�m��c) )���f�,ظc�M�os�i���E�����r��`!���7�j�f��-��1o��#9S��z�	��և�@�wC�>n�n��'�]9�ձ�f
��Y(��0�^m���r��q�\r:�~ST��޻%��5���5��6䨅�탢�l�T�P����.���4��a�`H�)���8�T�_`����V�㳺���H�u��� ��u@��Ji�^��S�w�ж��i�
��c�,�Bn�J���!�T1��J�Z�hd<�-�G��:����[��*�/�|�0�@$�L��N���N�ɰ�X�ˑ��V(ݏ洣���Z�! ��F �D����T��( ݮ؉8V�:N����~�ppY����3��ը���PY���Y2L�z��������=S��y�^����ː,�3�)����e�2�-���Dꅅ|�����U�@�V�ɑ�ȩ�ݭ����՛pa$��Re�MR�e�m��j�F�gr�=㻴��g(p]Y�e"�@C�?��w�[
���/&�n]l����~�Q�nY�T[5�!F�}��3(j_|U%N���]78��<����|[�]��֤��n�Qc>o$UpՈ�0�Q���fjpZQ3�ccw�I��<��3���A�ݥp��sZ�0k�k2�Xɖ$C��~3~_>7�ɸ�0l3�܆�n�w��eD0DJ&�I:��ץ�fϋZ�S�!l�~�ՓX
4�j�?��~<E�:�GI!M�n>�����	RWk��o�[�Z�b��7���L��'�+��#O.]�#�.��f������>зm>PZ��p���G�x$���'
I���O�Dɗ.���wO�����R���>r�z��N&$R��KMY�N�T�x7����"e6���;D�΍&T^kom!$�x���&��_����/�����v���-�� �{�|U��#�{�oغ'��d�8�I	�r+> ��b1Z{��Xt���Q�Su�l�HK"/H�{8R��&�p���!$���-��ܛ���`����IX���M�eF-�	�%�|��M�lYH �?h'k|���"�]�=�y���D�)�oF�}��c��T�;ܓcu 1g�5N#����q��z���%��8�������͢�B�ư���c�РC��������[��Ȩk���	�Ъ�~b�5����`� ����3�X�8�[�𒬞�	���q��l�qj�`-�����,�\Σ~����1R%(�~	,�%9
1$�I��Uڸ�?�� |��n�&�բw��)i�$���(| ���q��P����f�k����L2������B�i@"y@N(�w'�c��&(z�+�����uN��F�15.Dē����V[/�Wgct[��C�)�0.x:������Yj�����zW�ڰ9w����c�~�����O����!$_ۗx��O�a�j�fN�i+�<�{�
��J!%r���+�.�w�����f�vy��������d�:�/����N��U�H4D�~���y0�*4��o�T��Ͷ-j;�վ�M�� ���_>�RRc�p,u�Q�!b�pŘ�����[M�C��^ �񝊒u���T���3- B|�>�<]4��u"HlN��h�5&�"�G���b��w����0r�;���b��^�hh�|-Ee��.�����9*�_$R�*|�](��٩R0JIMlCԭ�;�ol��i�����sS3�`����S��$���~L�s�5��x���|wk�qj42jf�;�޻�FT�� ��Ƨ�_ԠdA�xeˤ7M��x�,�i+�~�ax�B�S����(��
����Ƨ擺�:	W�s�ﶻ�Ҡ��d��d���nj�I%�D���ފs؇�l	�𭋍!Q�7c:Z����iVB}qٮ�ͭ��M�Q���a �2�PmH3	⪕�I�V��8Ԑ�L��wz^�Fʉ�qD5���t�裍T7�����j[�Y��L�2�ތT_f�����Zd�����Ǆ���	P�z~�>h�����p,�~-�|A4��9�%���G���|̨r�V���_rg�ABG� =�P�^i�7��ض��B��a?����"�F;�p�T��W�4�x�\����1��1r"xۈ�Qj��6�$d߆���8)H>��B=�eE��1[��b��ЦO�X߈��e�X� !���ú�RU�X���E���Ub`ѡ�e���BO���Yһ�i����yg�*���Mq"[�a⊉�カ5�
w^Ьv�@A���������E�6̕"IG���l� EXR0��S�T)��l�G�(������n�˟@��^��m�M��� d����(m���q~��.r���-��� �>�M�2���\q4��.K%��ه��v:T�"�A~�,���ɓW�8�͙�뵅G>.�n��`_=�['m����~h�,�qMI�&�lh�i��iI!VF��!VY�j��Y'6'�%�k�{�s8b�E��=�'_-h�"��'	�'Gw^" 8�{[��Zo��c�M%+<���CF��,��̗�������=D?����H!�S�C��ҥ+���7
+.��"�����>^���D|��7��3�j�R�Ǔ0ǈ�rY���(��E�GL��ww��5Y���(C�>n���� �݉:l��7k�;��8q�RMI�aMx8��g_uL�Z�h�Q-�c�+1���� ���h���$¯��W�fpc��!����f�8\n������$�%��8e�83�a��"N��ލ�K-bc��b�Pj7�$��?��CQ��[K`I�+YJ�U=�c˲�gbo\�~�E��L�����/�_{u�*Ɏ�;X����Ie]�d���P�[�����!VAۑT�1���:�u}��,Jҽe�{�Ğp���r��S4�@��+o��D�1��Ӻ{�XG=Od;﮵"h�4�P�Fkp���y������GB萛��0Q�� +$D�#�>s�?L^`�v���ձ����-��8���{�%�����Gh�����O����2ư������"�Z���R�|>NU��c#h'þ>DN:�C*�\��۫_r�	1x�P0��Ii�����~V{���w=�o>)"]�#��J�m*�JlZ�4S�p�����4,E>�+���K*���_L[2�:D!�~���a�l%��l�Q~���M@[�D���(�^a-Y/�9| ��4�� [�j���v����0v�����\lr����4��@�]a���"E�ўy�s҅�[�Bȋ��>Y9U}�_֠	wV���\��q�b�f�ȶ������ۛ
]$Wo�34c��AKz 4��mG����aɑ���,�NJe����W<������T�fWv>��p �1��\s>�� ��/��[=�]�֢���.�!�Z�$5�ݬ�|Vq�n' �<)��
��&|?|[��X��Tf��fh�OFs���h"�0��s|2v;M��2l/�����4�c\�N@���a�w�$�ҡI����_CqS�%�����? �q�E�`< v�Ŵ?[��X�6����q粼A%�D���Al��h\G�{��_z�0�'��9T*��[4E���[��C[�hTa Q���1C�3���ZJ�5����c=�o�h��/�J奸{d݋*�(�7��%�z�X��[lC����u ��jQ4��U�{�]rq�q%��s���FU�1I�C��6���
~[�c����a9��?�{=�n���9.g�a����>o#iq���������_!�zt���t��	��!���UNC*�I��@_�a����� �pb9�sʯfj�F�\/չ=�go��X}Z���Iޖk��R��%a���a����VY;¡�0�ߟ"��(dLD��	K̦I��ڊ�6�Z2�X��q��#<�VءR7A�n�mDy����:����{C�=7iVF2��Ø���rQ`�]ݼ#��9��B;�c���nk�Mǀb.f�$�#ڥ�?�z�����pӳ^�����������G��^%TʨxSzղ��|�|��rBXT�h����A���=Ey`D���t��{@3�<n�1gE>B���	��`أ��[����	�ZN�>h��9ޒq���:=QJ>_�U*�v�Z3���g6X�@fR��F��Z�]��`sh��r)L�u��9�?��F���[9�p���׶H�?���^d�1 ~	y�ߎM��������T@�$\
�q8a���6K��rEE��m�ieq3�fBqSG��i��t���T��V5"����绾֒Q�g?E�&�eH�{C����y�� ���vt�/�'���+=������
һr�Vc��x��>��OO���IFu{�RO�d�3�o��i�џK0�߄|����!�����85��^�ټ����e�С��.!/�����n������=ìp�S>H#?)�������$pJ�	���o��C���nFO���T��pDg*��<nv��	�/7yX���BmPk���}��#{t��4ZF[gYE���ZϮf��_�T��O3;��:��R�RK@)���j���F���?�$����g�P�ޏ;U��tÁ����^�9��{W*���`&S;C��iI!S� �W����_�v&���ou�$��Ș�I:���y�%����7L��AŮ�R�Zp{t`���t��¾���W|���(�,
lIm̄k\-��y��#������ćp��$�U�8�/�s-{�Q�g�ȥð}��b�az<KBȍ��M��7������LK����tW�Q��n|-NI�KJ��ʹkoU�r����b1L��6H��IE.ꥹظ�YJ�3}���Z��2d�W�vE�����q� �V�ߨάM#1<��`Ѩ������,�Q/%g�>���_{�� 0��4�S v���͋��J�rb�9������)T������学��X�����!4���c�^̂���?ߪ[̓�M,F�*	&�3�	u�2�$zT�94���(E�(�y=υ�.��fٲ^��Y�!�|BL*N��ZT����~_\�AQ��}�t�o=sEx�Bk�V(��#J�n~������KC4C������d!�IU�!����-=l4�!�n���	N帪 �Y�ɢI�TmxG�Rת�!��R�xoXP�x4#Fz��P��Jxq��h�r�N�j�W�s5��d�qA���'Sk�]��u�	�@;����p�����"�k6��lO����U�T/�6#jy2P�"�	�jw�@���Y<褈�g��������gad��{�KgB�/;� �|C��GV��u�7v(�;��(y	��h_���=� �.A0%��3�c~�Lmm+9g��oU��ڎ]�h�)�N%w,�>U5��-��9�����[��7�� `�2��
±���2!��÷d�+��, ���{����l�6>�i:��� m9�ǸQ�^K쵕���8�˱���N��)~:)���v*tQZY��ˢ����V�Sy��7��y)�jţǾyycp�T&0E
=[+?5�P�L�x<o�2���JKa�����[Dj����/�٭�����^e��Kie��\�����o������j:}�UY'u\l��{����VqI/��X.�h1� �N��Թ-�Ue%��i�,2�5���I�"�'T�f�t���Y��-���
ϋ|U^��gۊ�2��dRa�����O����r��]��9_,�Q�[hj1�çx�0�.�w�Vo�s���� ��E��a)�
2�Y��1}�����!u�֕BC��u��������)u$�#��� �L�O��n�6���|.���u��_��_^:Ǥ��e|�A��S��k�.!>����Զ�f��x=���;�I���^�ǲx��}���x����8&`jW��`�w�}�JF��r"Nr���ψAn3�}W]>g���� ��6�� ��m�B��f�.t�ȍ(�m��"FR�x�]ʎ�0Efg�9~�ZZ<��wF�w_N�E���2����6 ���o����;2����]�܄����
˳�A�s�5ҝ5>������X�� �̓��X���a��GA�N���&_C��1�3W�%��[�]�M���9heL .9��Zx�-w��u-�k��;v�����@�%('��Ni*��@�FR��Z�	o��C�_wm��ۡ炄3<��#v���mo�Ծ��&��^Ɏ_I/m�$�q��]��󮗚��-V$Q�o���	�M$�4b�v=X+�Z>J^&���8��I,�)帠�?�r'&PZ���|4)��D��ҍ�ƒ;+tH��^�����ܖ�*M�pL�p�xW\�1skjr�':Ԏ����D���ݨ�A�"�m�;��s��d�*H��^K�-+��&<�]��+Q`$:���ȋ��x��$K��
!�=�Ô��j�|��.�;ewM�����=ɞ��0��?q73l��R�1����Kh�����u�y#�d�|��Ƙ�j���&��Eս9�:��#k��*���D����H��51/�Oq��g���!
�E�l��4��DR{6P��y�!\$�u������6�oX��v<k�^E�;�y�gk��z�b�u������&�\T�w�$�� XA$��,ĩ��g����0@t��}'�MN���G	:ƅ��Dk�nr�����~�SY�ÿH�Z���/JU��c68�?��_��nkÝ/8�3�_�����D�����ӓ1�҇��k��X2v\}����~n�{�3��~�ö_[��%�w�O���e)׀BV�b=|��Y�m�4��b���̐�L0�1�&x��>WѼV��a�������!�e���O�ʶ�q�U��d�V��N~Ts�-��P�|�J�.J!L�t��hH/�9<�c�Ee�^r�����cm�Ʉ-�T~@vN���
Ǣ��O��\���s��_l:�j�.��r+�i�o2hˁ*gԇ=��"��a��mK�M��<����Y���UF3�n
ŏ8���w%e�z� n�_u!F��e�
} [��+���v���ƪ�H��7`�j������	y�|�JS#��x"�9>�r��ޕ�@xc��Ĕƪg:��8��؊�bj��x �9
�eRr�u��NDuB_R��1��KV�fש���?�7��Ey��`c����^'7F�q�h4��QZ�`|T�xR7��>��&=#5V�z!�z�V�"�>JrH���l�@�"�n��H�2�$���/D9~}�J�������Yd��
�h�<!u s�Ϯ`7�{W�����5�ڈ��V��eBB��7̱�B��K����d»}��Ô�UhC���>�	��g�s�\�f�s#�J �/U�sp���|�	����l{ٳ���� �r�d/���[�Y��2��)���D}#O��\߱"̫�R��=Կ[��֑�*)a��V"�yz�{R�S��㦷k߭͢�7�������M�	�V5k7���#)~�r�ۧ�u��M*&A����M�����e2�ͷ�OMR떳�����yQ��ħ/���o|�:Y�*~�S�K�tH�����84,<�(�'WjLFژ����6��COL�Y��Y����@̠�w���m�g��7�=�A�m�;C�vr�4�$F�F�y���["�K�ϓ5�hk^k��<@�S����@OVx�0����D��&�.��.�Q��z<��H��B/]����� ��v]%�{�s����5T�>�z1��Z,�N�a�y:]grpk�6��O8�;�\�R]�0_��n�Қ�S�KC�E`�H��v����� �ϛ)�ld�	���6EOWAcBͪ��$u=(_Vs%B���-]��f5��.o=b۞�P�j��������ӛFn�K\�Y����p90�!�g��F*h��Ϸj��ʶ���>��q���⢤Z\��l���h��$h��n��z�S[1���L\�"�M׌0ׂ��Rc�����G�cf��o����eM�8�XRwh��/�+v�lQJ
�#�%!F�:��Z����G�@w���H��䫓�8uXC��zʝn֤��']g �6�	V~Ws\�E}�Z!�A#d����z噪6
�i�1)�م.ͻ�Mk���M�}�	���gS���H孓tq??��w�>�	�\��$���T�z��%�
�j@��4��e J��v�uf���<�y��~�3��Ԋ���M4�Ky��z�~oC2�+���+�*�h�&u�������s�PI�`Ƶ5j�M�ӷ-,�tR����;X'�oO7��O|Sxn
e�B���%v
z(W������C�X��$h�!��k׆,�p� n�a/sS���܊��b=��M}���>&.Q�I�q<����Y�~m�9@�pO�m�����f'��#Uf=@o��q3�1f{˸@��p��F�M����2����B��q�{�&i�p���W骡�#ڮ���Y!Ư�1�;�X� ���@���>��gt�6�\�_��0Q{���� �P �v�~{�hZ˺ߑ5���*2�G���g4�fl�`��`���j��V��c��F����y!*�6���5|?�=AX�I�6�Mq~0P><yt;�l���`�%�� ���U�$d ��I7�?�#��^w���IJ�\'�ϯu�ݭ�A�f�y�zn��L�ٱ6�=�B,�a�g�����Z!g����#o���w��u��sNK�.��f5y0㠧�_$��A��8Z0T|�4`��Y_k�`������w��Cf�`�]Jݲ��2���˜'�P�	!���dD"��?`E���6��
%�
�VRz�l�DnL��,��!6[8+td��/v-s\a���D�0�2	��{=V��f_��}���Z��W�t<�����X"�Pd1�T^�dՓJ�G�3ƌ+$��I���� ���f/�{��٬�gbX�3�'�|Q�X�Vgꌩ�t��u�h!���o��?�%��H�}��|�����h9b���e�.��F��o��s𚟃��e�g���S`3�z��^'��Wg�XXj�K��p�⠈p�Ƕ흨�t�x�H�v�\�ux��xZC��M�1�I(��Ue�H��FbkfN�wt$(�L�^�`Nֿ9��jW�}:%a�r�� 0��^j�y��tqX�	h�U�Xs�+���Z�vy�Z���H'�N�j��qE�v� ���Ƕ_|��R�ZJR��=��po'��i=� g^-���iz�Jp
5�� �z|�onGLT�-�ٴ��	wbHუM4К1)�W�z��~�Td�B�L�Z���[��[�0,��n[�#	k��׿�;���&
&��>�*o���6�aWL^9,�g㨿�ˁ� x۲_���MFm8��V�R�5����2\��j�:��Q�]V�Ht�?�S��̾x����+ۃ����u��Rnyo&axa�X�,�}e���U�H�gA�ʟy��R�h%�b=s�I�"��x�,W�-��e�h����	t7�;��*�9���[����������c� X騸Ւt��aB˳��+�K�h��M4d��Rz�(!O!�Ϟ_g�e�xU�q��ybtK��J)��� �C��w��~���i"��dr�e�.�;3�	X�g�V?���T��O<�;�}Ht[2�Vë*E���Ơ�
����y�l�����N��'��^���-G���R|��p�Qj�Z]t�+�whN����kT�@H���]?[܈K�����F cliv=��dI��V�?C@!@+��x���x�Nkg��.1�X���W�ň�7������|��ъ���m�&�۔J���?�=��V���D�,�B�Zy5�b�R� �4�s͇�AZ�R��O��g%���B���zC(�59�H1�r�~B�[}gj�j��\[�_�2�Ɍ�{��[���g��H�h�@ď�kz2h�b�jl��XU(��U�((a�R�������ï��p�~y�9�7X/��<�/�	^e�8�J`��-ϼ��y���nu��@milB]�G��Ъ;[0�e'�;�F�&�?�xJ��lz�y~s)a�R<�G̖@�1��4F#n,�G���`���:i�x�##�����Ż���{�C����=2��o:&���`������L��7�%!����Q�$�͕R��A)d�0#3F�w>�? ���I�'
��f\`hBrlmVȕ:7��1O�[->��H�ٶi̤��uњ���}�/�SCQ�mY��l2�Օɸ��4K6�87�H��"C�V��(�4X�]M���-���_g�<�&(�%@�>�fB��>�0r�ʣ�_�aaµ�VJR�����SQ��|�-��}���z���q�T��ɧ�҃��U�7~NE�dd6�d��q�w������J��Z����D+�XAK�j2��;����8��R��4HNh�x��9�����b�ʯD�xk�B8[A��$MS�в=4L�<����K�(������KH���l>��Dv�RI�aHu(��>�� �]����ULY�"�����,ġB��*�Z�&�����5����ժO���r�w�[��S��F3����$���_��PΠWd�h��r�Ԑ���x���#3�`<].��Z��&u{�e���Ć�>Gp$��QE @���4g�����/Hp��ahQ��ř�<����;��E�
�	�g���\�g
����1�ʟ��� ���p�_:��b�u񷤫S���]XG�g4����8��9�gF��\(3�����:<$���|.�=]y%�:ߨ��w�c�UI�f���7f��#7�u�����M]w
,`lB�����X�������V��h7r�Y㮯vO?��i�4�b�m0T�4U�������1#�	Ǩ6I,���,2���D8�A�g�D'@F4�ۢ8���Ah��Et�F�a����ZD� r���:� O1T4 �u�¡�ir�|��"+�L�����Q�f��;At�����0��	��r�yda2)ד3�mu�D���2<�����]�i~�=�E�8/gLl�X�/&��=.����5)E�\�.�֡O⹐٭i�I�l�Q�k<I6&���B���H����s�P~��]0�Tfe5������ٱ�=�x��MƘv0έ��P�W�i��F�ٵ=�H�:�^�ڳFa{y��SMT�.���\%M�|q�s��S�^�v�>�(i�@Ia���9C0�"�ˏm@�<KZ�S�D�-�a	[��yt���F>�`���*b/o��I	ـ��(�.)�6�i�T:���.>%�Z|eWOs���󲵟`VO�8px�F�݊�B����e�q���C��rc|e0�������}���W&B�i>{o#�\�j�����	 M� i_���p��]SK�?����8���l���sP���P�#m�t$�H�ˎ
y����:��8�o��gK���������VG�n$�w�k��QEx�����}o�U~�4�AJ����Q��|������k3�0��9���v��=�L��9�4��5�t��m�]�� �'nU�U��!��'�C#NgX�4���������:0:���\p)6t��|ܹG]�[~xNl�uj���eݚ�{�ū����l}�i饿���{�b���N��=�Uy���/��<�в�<g
=��3O
J
1�tj�NB��11ƗI������k��35�+���i
	[=B;��W�d|^��h
v�C��[M���[h]ֽ��h�y�U2Cn*B75D߱��&\;�_��fC����ߖ����f�s���� ��f��ky�6ln.:��znw���D>���K�-���l�D�$���jѻa?����<u���Q�0pG�hE�:������EA��5U���R��>���H�OZ��:���	!�p�#o���~�L
�]Y�}-����2��1��_9�~��^b��� ��Mg��uS|��Z��4Ү6��ӵ~�^�b%6YxM��K�_Mj�B�q-�*�u�i5-�mX��'#��BL_�ML���T�ǅ����qr�n6��5(�ѵ<�>x� e��K�-Z
�|�aF7,
�`<ҽ�y�|א�}��n6`[A���}�*(N$+`U���/���Q9绱��,j�$�[��n�_�!Pq��(�z=@�6�ײ٘�ެ���i��P������4=Ӎ)L\\,��-�5J�u�J��5�V#�M��Zr��y��,�!i�~�<���7F�� b�(�x�O�Y ����ɝB��4I�*	9墼���S���~��>8�]���'�%����� �eE�J�_��s��Nu�ڕ���-��oM�c�D�'E�G��f5��!�bK2�='�V]x��i����n���A�a���covʾ��z�>pV���J��v̱}S��Ξ>�H?����ަ!��M������E�Gd��b�R�V�Ν�O��è�Ʀ�2�b����T#}<"�Q���ʄF�G���٠�{.�<�_#}�����?���!j� ٩JPi�Řz&�k�,�3���չ�D�X�&��CjU�N��=��(���Z�%�/����� �cm��|=���IL>v��&צɡ����&7>�-'��b�}'eIj:U�������n[#�S揣@"?�u�qּ��t�ʍ�\��Ŕ�b����U}�K�����(eI�����ܗz��X�dJ��������]���h��mlĜ���fJAZ���3��w�}���H�ĄqTP��m$���﷬>=yS��L��q�q7 ��R�(Ӵ��$ά�u��`o�k�"&����͚U]ĞAi���B:���`�^d
h� 9�Th��N��X�;� �/����e�ը��"]�>���>W����p��,L����~#*	ď���U���+:^��2`�bf�~ڐ�W���)����4u+�H����)t9���) Q���y�kq��x��b�tu�}h�֗��Chnҗ���/c��OkpFlwj�������M���Xrߓz�Y���B+�����3ߔ�4Y��`m�۽y��ӏ6�"�1�j��x��=8��׶U㷑�xhQW}��+E�د�[���<B�8��!
��[癤���\7�����Zf�U��A�T^4�P�����b����������G��8��sv_�Ů-�+���C��1S�7[Ik��4_ N��X�>Y�!:)DI%��"�$�������]�i9���ts�-��:��Ӹae"L�i��b�
���*�_��kz �u�X�ϸ�ߋ?���~�ْ�u�Wh������ѥ�u�[��fF�}�.��T����'y�*��v���oД�U�pJ��n�d.RM m��x}q��w'3 ��o��b�u��4��̷f�Ve=æ�o���ais���3�!j,�����V�G��%An����P�ܩ���>֑�?�9���*��bݬ�.d.�eQD\��\f���������Up9(�˘��0���(A�S�-�Oo؋O�����<� (���V�x��5i�K�4f�����RLM$��SQ�`a��� ����ɍ�@̓;x��eP�|�<u9�$����~��^{M�Fߦ�n݌��{?��<ܣ'�CR�.Nؗ�k]�z�
m��Z�[��3mU���{��8�GoRnek��jTY$P]����Z�!�������6�'��p��|d�e�OyW哥j��R��͒���W��tF�A�u�O�%����d�4�\���!n��LqԤ�{�ZS<>N�L��M�.�֎�+9D���Sr�,������&�� �U�e�s��K��'@[�y�󼹞dt��1<%lg���3!���g� P'c��g<eK�xX�!&�7��)�(?D�8����Ss&�����@~���^T�<m��@;fz��a�w��u&�O��Ql�?�Ѯa�^����`K����+��*��l�5�Q-���磏4ǽj�>N	X���fj7�[!�^�Xl[Er`H�k�i�vn�1j_99�D�i�����-�W�[py�Ĥt�h�Q�L�p�̽��n�b�]�Ho��C�P���Ÿ��=�!����]�s��X!Eu?tt��Up�AEβ�� M= �ti��焄i$	1�q����M�t&"ߡ�E$ޘ- 'N�R8�5\���!Z�X��PxS�Wx��hXi������/��5���T2�J�z�{ h:H�unZ�	"�`���Xm���@Ɔ!4�ο����X���f��s�O�\^���q�d��@�KjQEc���?߰vs�*9NN��F������O>T��j��(]�{jd��LlN�pW�1�a�P|��I����wEu?�~
��!i0E���T�@Lyb�N��ζ��Ova����M�m���1��w{�o�\Gw6Q9{p��*��Y�Q{���i�eU�SN0�z��
(Ř-��m�uX�s�6^�LHr�Ӌ��ƀ\~{��G�������a\V���^?;�E�Q���r,X|�B�5�-&Б���GgV�����;G�;7ED�/-#��/���C��Z�Ѧ߈$B��g�����So<��p��#F���Qe����)-%Y/m��e��I�eH�x�jmB��ڟ���~��Aԃē��"իS�1�����ʲ�,ې�R
�ќ�ʰ�V"f۲|j9��Q0/v�tNqĄ�����R�;q��'nc���!:+�T�>,�k��c��M��$Y�w���\*Hgl�n@(F._~bD$�'�xO1_�ʵ�tH+��g�y��8�>���۾i�<pFS�*U`��.ԍ�#����x�Ӟl���+��N�@��'���kS��"�S�>��w�V�Kh��5S���WP[%TZ�A��$�+�9)�&Q�P����x)�;덠BZ������:�Pn�he�Fq(�խ`$���X�X�"�R��W�{S�#�z�yb��4p�qt�3i}}ƾ��u�ῳ���C��̣\}W��uY��H ڐ�B��g�BMD��-��6U�c�:���`,��.��Ā{N�SO3/6�52�L*����*wUJ����O�z;*��*�3NJ0���b݃�v��Ob� ��� WC&�䛨<����jW;2��kl~�1I�yP6$A��SA	��_�5��H�^%��Ƭ�2�#��by�1��$sʯ���%U�����{[�?c7�T'��~{<u�6{�s��@��(5>�����(��[߷�S��"i��K�{}a��Y3f>�I�(-L�ޔh,����7�
���N[F�<��7k�\C��|��@���vy�ҟ'6�ul���aª�\���b�m���U&�������=`�����.���_��쎓���73NZ��cI%z��V��Z�s�ymۉ|XC����)�߭�:�K>6>�S�M���d���TtƟ:��a�}��G�Dv����\�@�JGj�X�D���`(N}� [�P�v��_>��Iu[���A�k���%��H���ea%��r{#i]�4W +W�WY5i0t����$�^7c��2��h)\�
h��[�9��;\5����:^p���'@	
�� 6�Î�x.D��q,��I!�UR럾��	�Q��:^ Q���N�.i�����B>N��-!�-h49��T���1��5�؊A��g'��f�P�4דn:��I���O�&�'��s�4%m�5ů>q(�����\��6t~<�gԒ	1G��R�2�51*+�;S�t�sʰlm�ve��p��=��K³?�AF��I�C���H��h�,���Dܶ�(y��H��;�_��oe��+d��/9X�MMOX�c�:8��A2u,!�1>���?���9���C/lR�u�"�U��aTHl�dC�'ݔe�i>б���XX��k��:�:V����=D�����Vo�$����������*@��I�2�<�,Om<��z��ZTKbf�fԛI7�lt�ǜ�XF޷�m
F�?����1�w,��Ŷ"�����q�N`�J�����o��/�E��%�W�A�k�%�|$�ܳq�C=�.O3����S�5�~�Y:#��ӿ)�utsP�~,�l\*���*�)�6)�5�&��\X*���o0�_H�~N�����G@nժ�iB�@'H.�������ޡ��v��;a2y��0hl�l�-@��}W5�gK�X��E0�k��m"�\̴�>���dV���qK%�C�&b�]��"R*�%��e�`��}�����_�!8�x����^�v-p��cm����@u����6p�vR�3E7�D����?�MoM��b�mR��3i'_?ϵ��z�F��'�Ю�]Sd@m�ОM�Z6d���3Qq���7��D͢��,�u1��u�JiX2��
�@�J�;I���^��gˡMkEi1{����)L��	�6�r�������-Ml�/�b̲[���y�k���mI��jE�y�\��@��7P�6�+n�q�Hi�����(���j>��X�4zn��c�oT��(����O������]4���w��e�Z��δ Om!��k+_h@	m���rI��WY����J��Gw���%�y��	;���4�pUx����a�)S|��� ���`|�3&I�|L(�M�D�6���D�����B��i�%�c}�݂o�z*�f�V%�a����ݎ��q52��b�T4�H������c/�䂲�I��otuiގ�#�����Ӈ5�	b��۵��k�K���ȧr�^䈔��%��,Q��:�.���n6{�gOp�d�>O�=6#��]���}�E�V�������qb;�Ѽ�u.1D�!���`Tq߮�}�v�6ѿB�����A@"DV ��e�>C[�P�g|�)F�C���S�r�-*z��hI	�pPG�j(fhj���b�Z0ToT|��"Te��+��9���#���H@�����,DE�3����ו�܇*Rܿ�oǟ�E�؏���
��w�7�?�H�s.g����S�o�ͭ�K�g�:c$&�٭d���̝nh)ߢ�����5B.<`a����@�����S��"�FN��	���P��K���F� ��Y����y��}�����E�`�������t��	[�ȡ���,��a���Zd��F߇F��f�G���
�+�Iڂ�_h�A��V\fS���g�-�Q��Yyr����\�:�m��Mș_�8BE�Z�9�N���'F�7�?G��	>�;�7����<	M|�(�ah�xR֓ܝ� x����tv���ϭCT�M�T�T���v�K�^d��o��ϵ�`�k۸1�V)����[�Vu���6�,�'�S����PJ�_|?-w�e,�`��XSs�	l/P�E���!�cE��L�%|�6����$[�׌4u�6m* ��#���jfQUؓi�� 8�I�>�${�"��^08Z��1S�4��f��V��(��Y��i��mPI��j��ی����<X��.�������'4b�G=�}��ʣ��Qkd�Hc�����L)W2HȄ0�y�c��kx�bsŝ�vb��p��9<����ߑ����q��h��Y�%#Y�&���	vCT�M���&�y	�ޘ5���kh�Z��L~v���|v��N��{���%�h�d�j
Sm?6��8����c�_o�����̀~| �S���-������D��C���j�Lj��� �|8#(4��-�� Y{eJҦޞz�F��!�5��]��P�Zy�!@��cy��������(n�<��9�oj�|0R���g㙁�'���(Fk�Eu�طwj�&�թ�] ����F���
�P���s�n�0cPӰ[R�J2�eIh�%����1���5?+��;	��8i-R'�S���E�D�i��Vc�n违ӓ2V�)��3��(�a�A�ӕ�(�}Z�,�6I�m�Ѹ��?�Pt&C�&����k��Gu��R�`B.C�/��j~��V&ǈ���.������<[&W����.�V��;��?����o�gB^Y����j?����
N�904s���H�w�o�;��ù�sp�9)�&��D)�
��d��p���'�4�e/[�Z$�[�"��� 熤G����o��Ò�7����oEm�{T��٭L�j��V��ޚ0��R׻x]�"}�$)�݂K0���#��M�&��v�T+XRJ��Y��Gg�����G���ݧ�M2���U�zet�^"�����	ٙ�a��#Ti��>!n/��H�@�EH+���@=���E��)n~�p��[�"E����\ohw4;fzU�F�>�b�**�1�HW��j"�HɁ�Qd;�����Xd�Ã�#J�H�Ǆ�دcWe
�X�I�{���A��TQ^B��.^vX.� ;��uox(�S�/*5��۔��0#�N�KH�{Jަ	��a3�8Y�(%�*D�7��TzV�C<^�-I�
�y���lcj�J.R��5嚁��x6��R��^3!߽�ȣLy��;��썱��Iт?]ӗ�*�)�kv�`��c%�+�g�ֿ�OzZ�Ű4͘���g�n"��"�?�p|Q)��-�g�m�.�I�s�}��{7�U�@(��CH0����I�,L�8|�� Q2E�T#�w�<�I�eS�c����=C�݁M���ꗸ�"( &f#w+L ��bm4��$@@�fKVz����:�4�s�	鳅,m=�K��[�n�:�p4��Ru4���
�!�5�^?�'��	 <O�?3�r;ӥ������?F�π{�ˣ�����5��Y(������\�~�RCT	ޔ>��(�M?��X���;7Pƫz��J�`�1-�3�2q�;K�㟽����xU���뜵|�D���(*�CO!�jO��~ok�/1�+�%�/�������&��X���\Eb��J����Ԥn��5#1�*7	�_�����{)�[,[t 	#�u����^P�/����ӊ��A�>�	�ݏ?����_0$���ʽ&�T��W-�f�H�ݏI����������I��AH�a�
�ˌo�����Q�yn��T9W݆w� ��.��r��Ĺi��<
u<� ��s^���q�N�nˬ?����љj����SЁ�4kL<-Y/�+C6���h1T�+JB��CҮ0x^�O�aҮtN�.��9���:�*VZ����-����Y7דX	�N���8���I�
�F��I��责X�3,��.����,H�愯ro1��(��6u�%诵��UD��Y��1�!� �w�x�Tԛ���ͽ�h!� :�b�WT����e}Z���v"�����b��O�i~����{���b��&����!���3Ӓ���X ��|TL.�s��z�'z$�s����n�\^��M�Z������v*a�8-L��NZ �>_�#�V���k��~V�hЉ�T��N��A+���
��>�6�צbq ���}�Ҍ�k���9�S�c��x�K4�'�+��?�y2��5/R�Y���X�B+TWA�~�]����ŗ���4l�e��U\o��������2�>��lJ�!>1^�������)��M� U�O~�,#992�����:%�ܮtx�pm���]��L�vI���4��x��TܰTb��6�Q�g�Y����	[b�jsPMa�s0\4���;*�W	.yW��P�m�N �iϜ�42�9W\���lI,��BZc��%,������6,�R�5���y��h"Y��E<��|�?�d)6��'�F�~/E�d�����d�Ja�{����5&I���T��$1Xtn}��l���������I�`���Jdu�؅|z�I�AZ�z����~�f(���#�=�/-;R�U8~�5ZM�6CV����"spB��H�|�?�mK߄��ѥa4�Y�J���ư�Q�_�=��,� ��""U+V��F8���r�ki���,M��A�jg;���e��q�$���D暼O��|�ط�Vh5:��/up�Fڤp&�#G�g\�q����U8���'��i��d��谴�Bhq�~����(	�i�B C�O}��������>El/^�^�Е�ԪGbLP�s��[�"�*��SIhe��pj�\�t*f�?����e?A��2�z�R�%H��$B\��t ��g)�cۄHѰ����&5{̹P�i������J{�X3�x2.f0q�D��0��p�vJk$�j\��.̆<D�pI���
�.�؈�5��B���:��*a�0�M�)(�U��T��̗�⚥�g���z�]�<��J���R+���x�%rM�l1���@���~��5��_�/�`K��2TL0�ɞ�*�*%�2i���*�Ѐ��PPm:"f^>~���@0�b0<5���>�~秀	:�����'�A�P���g�V���C�c��/ ���IlN�mq�,�)ѯ&nK䟉�G�Š����az����ڮ_�H�ѡ������{�ꈉ#�Ҍ�u��!,H7K˄;K��0���u�y��a�D��Y2M Ս�,~}�ޠ�D��m-���V��+!��:B��ұt"�pPG�b� �cX*��ڥ�>D>(Crr�g�lA�u����ޙ��h�B�BF�A� 9J�6yS���q�1�� �i`�M�
��nAM�KI�	�9"rG�*��ĥY��e:�����x{����҅){�Cy����tKZV��i�����O����y�}��+�tT�r.㐷�{��̚cx����Q9g�"�x&��<����w<3� �=�k������ᶈVYw�>��h|������B�h�t�_j���m��Jˢ?�&K��SF}�n*�=u������q�ٳ(s瞼nIId��(vX���SP�D�t�lq�����Ww��6P:���m!ںh����H����<�?� x�M<��-EK^y�T���W��Kd1���SP+�z�UQ|�	�0��|�J'�n���Z�+� 	MP6�>t\Í���]BI �5�����r�d��\P�-���q�c9`���/���4��@�&^Q�6��$w��-�4���_igt ,��5VO=�|�&�'�����@Y�Ѳ��Q���ס�����а���	���4; [�� �?�֛�	�*�#"Ğ(xP�N!��05�䡀)[>'��	��U���D��&�(۱Ԙ�?�o@!Z��υ�s䈲.¼j��t�)	���7Ɏ�/k �b?�t����w7�{ �A:5�/m��9�B�u;լ�������7���������;�݈o�ėh�z)vD˩�@ '&m<կ:6����~>YX���Da	{9�����+��]��͔��	�7 Q��O���N�B���l�޾Y�s��;�<�s�$�&~�@8U\*����>E_ �f����O������R&A���`D��?�oB��#�M��W�"/=r�3%��/ػ�a�#L�֎w���,ي�����n���n��<��Ur�GI�q�Q���Z�T^8�T!r���uf] �@�dk8���/���Ơ+�:Ȟ����6'��O��2��в�]�]���=�Ge*�;-	Et-"��2�_v+=��}y¥�
z���hK%	M�v�M߃I"]�=.)},���)l<P��n��M�-����b
�I7����7lU�t�d�Р��ԑȟ�dpU�������]�ͦC�&㛼��w������S"b�X��\0��TX� L�l��}*�?@�rS5�;�x��ɍ�6��xֶR�p&��z,,���g��?0�Ld�e�]	�|ҟ^i��!��M�N]���`�Ez����i�s
l8
�j�-��Q�\-� rlx�$��ԃ���Ja������%`2����T��$P6W��c����Y1���$3ǋ�l�pϓDh���K0��}�%͞	��C}0���͐�P���nq���H���b��l�����X��H6?�+�"H��ݺ՚�e�Ҝ���%J�9���<Q��Ǯ]Ts�
�F|wfs=[���Aq�P�r�H\G>*@�sɁR��h�2ȨG�tL��J�5��
��w	˞�7�j��d�������p���1�2'E̾��r�>��z�Gcl�$�	x9�bP���y�qu+�ZɐQ��L��Ho6��dՀW�CJwjs������?������Z�kl�7��8���)h�V=mS��i�W31�yk��!]v����ubn*�F?h��L�0=�6��H�,O�N������.Զ��O{6��]��2��]�5F`�`�Fʡ�A^�2�+h?Ĭ8jiG�W�0����l��bJ�H�q���.��t��L��L�����2��q������o!v��@�	.j%�w(�r�jc���ӣ��lc�d~�;��r
�^����6��Np���n��W�זև�-r[}р܅v_�,+y�LįML�7��<�����𯿽Z�\_S��f(��vs)�v�zܐ?��~=u�t:㷩EU�l̀�eKA��^ݞ�@o`��.F#�u�,_ � �r$��}ͮ��q	��j���?g�bx�8�{ kp�C���.�6��PN��5x���Sb��.W;��X�^����q�8��֏K6��Չ�ٻ��5t<�C���a.D����<�'�Yz���D�xb<%D��zS�!���+�P���B�LU��ѓ<�}���`\v4H$��!�|!��a�*����>�|�n�\���5�;��W-��H�	^D�>` �|�(�|��������\�63���Ht�v.R¢c�\E%���s@b��9�}]'p�G���*�ζ��O	L(������|w�Mo��eU��`{�>��k����b�k-�sy�d#�틕�7|�iC3(k�k����B9� q)o��C"�Rs�/��	����_�̕�6eY�F��ԥ+����i�L��{x����p�&G��21ũ1k��T�k�!�(d6�Pd���������Q�('R�=�5נ��,P-N���>��uy4�	]��X�.���h(k��v�jXS��r�=���� ��9���5C�О�8�u�ϓ�۵�=�8c���j^�������N�g�[M_ �0U�7Uq��r����3rv��Lz���/W+(��h�|�6]��
cA����u���aU���b�߇u��sqV/��+�@��mܳ�ÝGh�p(�,�Z#c^n,�{����.�7�I�����k�1#��J����a���l����`��I��v�N��ԍ�;:F��0�S�u���ȯ��^���c-|�3�AO�Y��,�G�D;��� �l�# 6�H�w3À�dr"���0��"�)yk���?u����_a�ۂ�gN�^&�>��*� ���eWG�o��%j�Ђ�Nܖ��H���L�leǥp �]�aКy�hL�x_5�Ýa�d�H.fb)O-/�H��w�x�?��໨Cl�IUMBº���G��o������Z�g<1�-�k̪���3r�K�N�����/[�]��X���/���J�C-�@	�e�Z�l��B�#<\�!4v9E)�#�E�/�nr@�~��u}�&��y���e�V:N���>wNb
[	�l��l���h�᫪d�j!��0vNn��ni"�̄G@4��@�3�e�W��W�
��V�O���`�D�k3��/�9�c�� �$�����P�	�1l�&|
d�Ϊ��f�������E��n#�Q���>=�Ey� �{Ҍtӽ�*Y�I9z;U}���68���r��E]
)I����bx�M �:ݔta0�6�?��[���#t�a�X��L�'�b|�83��	���:���;��"�{f&O�)�m�6�����[k���W[6C�����l�r�"�����z�w�J�1�ƛz���}�I9ӕk��2,]48d���|6���UJLT����rˢ{��vk\}��6"�V���^���|��+\0�&��n���}G���-{�<c"���
9��]k��D���Z���]C�N���簛��alW��H�O���E���H��Vy_�5�	N�ͫ�|q���m�p:3�v)v
��IH��d ����0�.�/mK&���g�6ΈB8t�+ˠ�����Z�^&��9���W]7�u��ӫ�Qm�B�����v(�8�;�p�[���H*�XĽ�B�#��:K���K+C&�%�W��-���Ke��0�j��=�~�ŧ~�yv��*��wYt���%��Đ�2"9�~w�ă�`��h��Ҿ��0l�Ul���ط�D��ܺS"ȷOni���	l��V�|��tB��ۗ��`1
������������+�ϧ�� ��7� �8�ɏ��\yEIgy�����,�Ev)×����ut�r�K0X�Q3��b�Tٛ�>�d�C�;� &	AÊ�`l�U7�h�/#B]
��D��<�e	m�vo�@��t�H\�8���V��*υ��Ѻ"�!��Y����R7\��4ʪܴ�����!��ͷ��)��Xf4�*&��l9��|��p+R�Ӕ��g����EZEY	9�2-�-���n��X�kY$у��8y�����,m<۳T��4��|�w0* iӰ�a(��W�JbH���坰K�&��D{��z`�ڪ�����N>9i\5��ݐ�
�� ��:��Q��*L"��֯�5�Q����Z�3�s��?��]�P�Y���������ϙ���9>@������*�g�M�ˣ`��DhO�����1n4{k����$��׃^��?r���x�>;�	�}׷�>1��/�YtF�y���N|?�G���y�&�Q�xITb����O�7*R�8�
"<�|Q���-^�p�Q2�\�ި�9��|j%�g�0�6�Vx�d�*|6H���Kƫ�PٓЖc�D�F�c��҇�Yp��w���?����׊LZ�Y���]��V� *�q�Ÿ��C]&�[\���Q*B�Z��g�cr�� BƘ�������L;Ks�~�g"ʘ��"� ��m����_���?�����lz�*PdL��%�/�0�u��x�^ ��t&�/I�3K3��L�E�9u�:��-����S|��q�v�ݳGtc�.F
��5��%/j���]�D I&$mdU���̨�<�{,�)Lv���[rrF-a~����%jr���X��KC�4%l��wYS_�p�
ܿ�B��_��邞'�8V��>�b:t9�j8������c�9U������fĮ^��n��|�_0���3�����)P�_
��M�Ƌz)e�Dmv�;�%{u	%��{���}D���l`j��f���N�f3��TАz�=���%���ĘF���D
�$E��s��&�И+|�g��	 ��0 T����)�h2�b�Qul���N��˞
�z=-��#�[�E���z������]^J�Lc�=�|�;Im�"��������[���a��|7�07��؟�A6�c������2���,�"�6�n>C��'�]�	%��hԵ`��������u��Px��6�p>/,�J����Uʞ2r���o��e�Z��}{3�[��:���o�Xy+��q���u`��:�C���(�u�〈Iw�{x�Hh���<�����C��bz\;*R��0ai�^m~
�KةdU��y���Y��6ʀ���fu�9 ���Vl���?���������H~����"�= �Rm�/��vǐ���wֹ��!F���ML�H�Q���V݌��g)���"����V���s���=[4YK�2����V��3�����|�m��a-��K-w���~�� In���{m�W_w�h�}��G�<����%��`X%kM~N��SSK����x�-uj��%;J�>�@.�Z�:K|��L�W�ص�V�b��PJL���l�u��	D|���8�<5��|i�գ����éR(g��u�6�͛�����s&�O�Rp4���L\�#�Ht�����~��i�z��q8s@���͆
���� ɏ�����b�|��yc�������x�Bb����Q�c�"|Qkx��vh���
K�fC�tS+��w9�Cv�=��2+�ʜ���?R�5��,���Y�}����8I3LD���97ҥ��;a������\	/>_���W�u^=�����b�JJ7`Q��Z0�J�f}�#nlz���(�e�Qo�V�#�����<�o]���9O/�K'ALK&O{�*�{���r��{�+b�2��q�et�)(�J%M_^�2���ьa�T�QF��Q�|��`*�ߑ��`�r@��%8�4b�
<�P����z��O�@i���;�����Zͫg��EիHg	m�?�0�W�#��|؛��?s��O>�s����E�U�t8r�O��h^%�9 ���I�}֚�3jMz�Y38IP]B�������Ȱ�p�ң|�g5��^�:�H�t�35r�5gY�F�(�p�&ܵ5J2��XK�.}B����S�Ms;gn1A�6���.A��Q1S���`l��Ω��JD�ivy�\u7�u���mnG���"��ua~�ۍ7�|Q�\�&Bc�W���TdW��t�,gנ��6s:�8ܑ�n���M���<DRFޫ�H��7�� 4�۪hX�I�,&�֮Y����2� �*���U�cM\"�(]��עjj�m�t�_W��ftf�3�j��W���%EC"��1����cO��!>RlP��v����H�_uO��"����I�g�&W��h6��� �+W�����1o��Ç��Ҩ:�w�9 �XL��速ئ!�W���Ș�+W����sR�拊(Աs�h�|��8���	�z7@IE��3}�m?#"������*�`h��0�8^[�f�:޾=�˰yD�:�>|�mu�(�2`ݯ[�{��Wr�������a>M�������A�ͦ��u���"�<��R�M<� 9;w�C_��k�������i�ڨ[�R��,=��16T�㕍^R���h���%_�\$��!?<Za~�*�:�?g����9w�L-�w7�KRrܽ)>��2��w_� Hk��[C;;&�ޡ¶���֦�gh*��ϑ϶�vN�G�W�t�Qj�r���C�DI5VI �O���C3����E�P}�ĭ�l{ߢ�.F�
�pC��<�����[5Ƒ��g�3[r'�x�#P�F�\2U�]+s���z�W{�b�:�90c5eMcA5v���#�'�k��ιJ�B�L�ٹ�I:�H]���犿��IzF>?���6 ?d����4y*�5|.8�"�5�������#�i0��g��-���*��M��>��XS����0B��B����Q��ֻ�]f��R8��nf�x��ؑ�����]��Zr�s�����T�����/�䥀��/�CЯ�6�$]��Bv����)�L��|�"����_�?�=҆�Dң��G�<�L�HD��I���}��u[�߻`����Ӣ�h������ip�b�g��׳� �lԻә�'�������D��~��ZU������Ԉ�f���94�G��swN��w1���}�Mq��Ө;�ޯ��Ks�5K��Ԥ8+��o�8kZ�R��0�/u-�A�~�#�0��R&��i(<�O3�;.�:,�+�-b���r�CkZ�����o�(�Z�~7�k��zuK���Ѹ`��s"8��?��L?��W�)�V[��1�DGe���Z�{2����^��2��`q�zz���C<��CGiЉ���8��P�3v��S���;X�ߺ�s-��e#hFo�t~�S��8�q�noa����d��+o��c�y m���;H�iVh�l]P}ߘC=��; 3in��K��"�K�Z3H��2|SW�����*��nm�B��Й���>N���S��Lݏ9�0Ȳ�pK�s�b��M�����F�m�P5�A��֚�W������1-"�{���G�9��W��l�1�'��DN�Ɛ'�k�K��31�?36,�,�I?�Q�3�r��S��>���^;l���fyX�f�u�s��R��ZA����Wk#�%�˅i,��{�B�ƈ}��� ��i9�*�G	(��|olSOph�>ӛL����Zc���]
���O�(Ni�oCj� �&N��/�̾���)ڷ]�f/��c\e�c���ԇ@Wk^�<��F:����j��EԽ���zҲ��-�m�r�4Aojg�zk���J��;��E9:ϡO�rdչC���ƶv"Zjw���ly6���ygJ��wW�����z}�	z~����`�KD�fL��ILnh)L�)�A��J�g��q�;�Ġͱ��f OH�N�6=�9�����A�-�Hc�,�`�7���#�$�gL[����	S��*��U��_��I��9���Sp�[�`}�&�<�~38����@�@`F���+�u�%��i�J`v=�8��j,i�LC*��HEq�8����A�S�7��,2��za����Y�g&:�lkD�Xp�b��1�_]w�ǝ��@I8���-��0���!�Y�Yӝ�*�'ô���&�"r�72�^9Zڃg$�D3'ZB�ʅ��1�������2��� x{~��C<-RM���j$���g7��aZ������Q,a3'�����V�(Oh�L���M�yMJ��>��Zc�u�Z2<⿞�4�A�����}��r��pM����q3=���mi$��ek<�����;���l����0�*m�����o)U�Ƕ��>?�aj6]��psiL�F��l06�� ��"�R(��������Z���Ä�ӥ^ �(S|�cT�ˀ1�ϧ�~ʹ�Q�Z,SҞ�:%�b8��~��9T��n��D�S?C �Hl�JO[�X_@�J�G��_<з��&�r; �&;�/?�°o��d���dʳd��� ��n�[�/c4��s�Fe�.wnNҽ��n챨wy��>G����ߚ�v�����{�Y�o\Q��F2'Lֶos�.c �3��2ef���m��(EB��'��d��0��NԂo!�NѾ1^�#ׄd��ӯ����x�n*��r�qrBh��Q�t����E�j7f[��0\
��ͭ��_G+���r����r<�Y`�}���t�{2�SY���iԶ�X&.x����=O��MV1e2~� w�NQ��0"Ǹ���?�_����5�}	��=�~���C;��>o.��"�'���ԚF=�$.q{�m�Yc{a{$'>]a,�)��GM�*��#�>|<��7��#�sEq��D� `�zI�T��.�� C�NY��!h
�����yRը�6��|p�9�u���4�S�����S3�|��V��SB3%2=q#A��=o֐Ҵ�|7�:Cs�S�5�����^Y���A`�E�k���r�
BT�&�?��������o���{�<T�a���, [TRlf��i�B.Z�d6�ȅh�,c���ikni�;��a'���2��ӱ�P��8Z~v���@F�b� ��!���!����FX��X�����=��Kq\��M��Vx�Y�X+�B{j�sk��%	�ʃE��Y'� DY�LX8�]�82J.H�+�.���H��e���Gq�.�p�y�<
��5V�X'+��,��q�<������Wѣ�t�RQ�d}��Mo�E�,����6�ӟR>���!��m���m��S�2z(�M���#º��
#�px1�Cۥ�xϣ�5�J;����3�9�;��Jʈ��s&�����=��P�-2�W��Tgu�s]�[�Ht������4��3x�7��d�#�dܾ�yи�,��P8���XV9��Z���lfKm}ξFܶh��$�k_�#��o���1�[��:ZB�����������VG"ץ_a�c�� <��@cl,�!M�c��0�:���_�U�?WP~��G  ��yjbB=�5c��0\�\l��D�$��Cm����7��}M�+�(��1�~�[$o MU�BX�12l6$�*�u�]�L�A��I�_��7����o�E]��/��FJ����0{��"�Ԇ�r!̴�үp�T�x�6k��C���Ԋ��C?-�8Ņډt9��5�t�=(�\�N�O�
��f\���2M^ ��z��?Vt�ޮ�U�ۭH��x�cw�� ������qI(�}����Yt.�"����ޙ��$X��WJr��H�I��3��N!��`���v��Ե=)�* �M���j�D ���W(��*P�V	M$�ս$A����D:��-��dH�Agp�zG�3�H�C:�%��}wY���|R����PE���4���ݞ{gK���D���T�KNk�9��5S+�ڙ����#=���0�-G�H�?g��*�d�P��n�ܨ�*J��9%4�^u���o�J�%�@U�/r,h_��P��F��V�q�Vd@�q�4c�v�cMK�Q|�_�Br*U�d(�]�L7nRko�H"	��/�A� "�+<� \�$s]�C��-ǅ�r�d:ų��D����s�"��d��Ry6�[���C$�II�[Ĩ+��Q�n�������{n�xv�A�9��)�����+����Cj���a��tGݳح�q��=���C[������R_���7�NJ�,��)G�5Ǔ����hBC��i�3J�
u޹]�l�ꩦ-Ѻd�JY#]��~i/	xG�G�8�7ZLI�Y-�F�ѻ���tL5�o�����@W���̇o��� � /0T�)0��6<�j٠먓onJ��-/r��i	v��'��p3��:�X�B ם�$@.�c�fdળ�MI�6O�$`��H�u�MlY�BҴ	�!K��ㆽ�ϭ�E��� �`v����Lvѿ��dƸ0�W���H�I[ԏ�%{/��R�������C
D�_�HeaۣH�t!�!���Hu��m���sLd��"Y�<g��S��'~KA�y�{,�X:V�I��
�JX@K�W �&�P/pM�DU@x3śh38��hR�%Q���`�u�E,�@���-���ˏM��Xk/�Q����8�r���@�^E�V4)V��f�����j#3~�^���17���E����-O5�kF�Vy��mI��67�������\�B�M���'�����5��p��B���x�A��L�}��ŅF���݆W�]���>��P�YD\�8|�>1Pb\H�����A�sҷ��j�;l0鰖�������ŌG����1�w����
���\�2� �f����fǮ�S��k;x�(wA]���߳����H :�˹�mV��HZ.��_�"q,Ls�	�������N:��*�Ó���P�ð�tc������1�3=�/�E��+;pfE�"Ǎ�Įb8�3�&k�q��b�S�t�E�M�t����
��U���b=�Ж�δ�EXBW{r� �j���y����
�	��I�{�#���@K*xR*�r��q�Y?��j�j�ކ�h�S㰁v*ch,�k�Ѥ4<E 06�3�8$� "q!ea�ek��>���׵�ɜ?.�x�.,w����1O|x�q�p�'q#B`i�4�Уw�+���)���O����<����q�Zi�8���z�|ԨC���Iy/�����D�>`�g�����$�V�i�0����(�d�Y�&*�}-��� �d�-�_dx~so��Y���`2l.��4ı�k��Y�r�s嚅0� rQ́���&qy�Aҝ��@(��j�f�ZN-�_�v�c*<�6� WοJ>\�]�ɝ��VFӐ�a��jnd9��z
�!��:������ezH�尿�ߡ�`��e��(��6K��Ȓ9v��Y�
�Mj��`6�<��y��	0d7�� ����1h�N�	�]�qF�����ګ�MeҖ/�e��e�˾�3e.���R�m����"n�h{q�K�K,�¡h)X�5����~mE���I�O��m.�1�u�c��nDY^<v��Q-ąV�����{Ҳ�;��k&�X�#"�/a�4у��@�	��<=1I>N>'��4l-�r �҅���o#7��w[����B7��Z���))o�z�"}�)�:���E�n�z~��5y��o��`����� �����Z�wk���f<���x�C�Э�?t����K�S��o�����n�X��X���5U|����h����yU��ͬ�p�̊Xs�\�96X���z�b�@���1�9�}�
��Y�r{b}(�m5�/(	�I�C��Yf���e��!�o���.@]�v�q�M�:\����̰�('if�'��g�/��>El���N^��1�����&����w��4_0")�|Fuc���&{ �>�4dv�h*ύ�\�����b/M���y�Yj������9��~K*+*4�c]]Bʱ]��O�Q����y'M;���P�8���H������Hq�o��==�X�g`r;�M,l�	;7 1W:NT� BY9f��U�C���Ǯ�*�C�V2��BI�Z�L�MBz-���D��@��S��p����j8l�G\W�ܿU���W���{j��-�IlJ��xû-���L�о��6AN���J�����t���!1qhc���i�����~�z/Z�lK3��I^�z�><���A�
[��K�7���
��Ȏ��/3���
���G��YeAˆ�n~C��#ؗ=)r�%��Y�Ũo�%rR�T���݈9��/#�A)u��mV�so�U��3-�ۺ�;�ً�a1��8 ��bػ07�����p��Wn �}����o������Tק62(��t�#c�}5��ߪ�X���ͳz��3��5�q��9X��CW���N!�Dr���ٻ}�L�x_w|��Y�Z�(��9��>lkDQ�ptߞl3#�(�+	�zX{�����G���W>H���y�SK�|�G�d8� %� P��<��l�]�<s��ŀl��P;���~��4����'��_ PϜ�S�@T�A��fVI̮���a8�"m��;��+��.��a�3._5���,�J�z��P��V�����Ik,�GNt}ہ���)�H���֯3Z�4����Ú'M��Hē�>�5��6�NK���#�pM�j=��|���>�剕��Q�<���5$���򟓸���O�� ;�u�,<Z�oM�<0�V�"�͹~0ox�,0�͝�Ug�	K�!z�'���e�$��N�n"�h�cp]� �mٮ���I�B� -�?]A�N�H��[�Сg�	�e�i"��4[����տF�����l��ķ����n���$������;CN�S���E��N��jf�\ٯ�dF����j�v7Z�e�<�ILn��H{zҙ��n�wwj����jj^7��P�}ݦ���+�5P�L�`v���#�^��jު��lj���V腦1/B*�C)V�wk���*�1'>�ri^�j���E2R���+�{��Q:���yf;�|h�0���_������N����ꡂ,�VZwl>on"�
�m�����n��%p����T_B����X%Mͳ�o?$^��3 �3��z�z-���D�ZX��v�c`�1+�v�<}��x�5�n4��Pr�>8��G�v�jY�;���n�dT���Ek��<<�����ʛ�_[�j�:��|���L���l8���A��y��Xݘ];�H;�s)��G#۩�*趃[��湂�l�^����F
��#)d,�p�R�]n��t�J�G��x����X��f�ع
9��O�Sb�G�{z�AO�T��o���N�M�3���u;��~!�����K!K�Q��I�����۠��*ue⚳O�b�xIJ���n\�#E�+��ם���ia����	o]���-��ӗC�2���[���P���s�O��u�S���y�"���#��g�&C#�����]VÏ��S���# ��9�s/��hԮ�w��V����8:�i��K!�"	sl����,9��~)� ��2�x��V��'F~��E+w�1tV�林�t`�xx�n0\{�l�L�M\7;�<�]���8�31P_��)�[���6PF_|쿨<6�<���I<z����/�@�ε�dt�n��7TAJ辪�~n��0����"C��xo����:O(F���w�����Hp'�
cL�=��`��3�C���F:Bc���F����da�sɈY�}��O����]�Ǉ��3��`��X��U�"Y��j{���3 h.�����V����
��%�Z�ЛO��k�&0�|EF�9�;��S����3����������0��b��k)Ô�Y�F�Wzs��0F����.�LO�`o��ѵA��aWx")���t�?5.���4�Zq��5w�"��(:����g����)U`Ⱥ�eh�%�Q���H.A}��&��~���e����i�o��:��9)c�C�7�5�=���V���7$i_W��d?:(��?*�-�`c6J�ץ��ee���.7����S��;͏��(v'lJ����ެ0O��t[�8�>��[B��*[��U`��ئ�rnU�R������I��UZ?Խܑ]��{��/�.'<W �����H��يĐð�ܟu_Q�����D�n}Q"����3�����M5���7t������)�D�	Kh����.k��G����X�i�#p~�v�rԿzB$t�!����Y�aA He�z;�A:�L��Jk8)�3_^���<p�Sku+�޾�&7�{P���W�E��ٴw�����Y������c�����\E,Ȏ1|��<t�Kt>�t��[!���{Кڐ;�QL68Z�E���z�a�/Q~���c��`�H�l?jN]�����5f��J�%r��1�o��L��B�^q�V8�O`x��З�4سy�%�VAzY��[�I�A\�PT�Ԩ)d��o�dj�v֦��@z�D=�*璟����X�s�83̗;uvo����zAe�n�ٯ3ڲP��* ~�A���`�:��9��D\9t���q�L( �ӖM4d>��Y!c�@���Z�DV`6�^m�~�>T��N��q�����5 o���n��kkv��b���E)4$i3���~�hvO%c��l:��E��C�CpI+X��Z�,Hr���8H ޚ~ƠP�*;�]J�X��
ҟ����@*ʲ�^\"������M�~Ț0
(�=�Q���i>^�P��Z<��%���.ZU SQ�]�M�S�à�'Y�(��5"H�~��AK�����sn��F�KeB0+�51&�=֍�#3�8��*=O��r��*�9�7:蟍��H��L��Cx�iس��Sݵ=�Ť�H����.tY���A�)��3� 3*L:�G�W�DrLdU\���bsy,�+:L9!GA"rQ�w��;[��!�{�t����w`!�2��<oܟ��4�f;u�+��̾����B�X�B�|�(�+c���I^o�k���ʌ��A}�$3m�$���yK���C�Jt�WR���Y��F
��"qDz�'A!k�^����$o�>�i�S��r�'����%���z0��Q�h���CI�+�Y颔X�-GD� ��<)S�!Ա��g�{u�U�*�{�i�����t0n�����4�9F�s��@�8��p��`��n�1���|�K�P����aib���wo��E��g��nχ���]{�|�~���(�[�G\�K���֋\c�t��6��ܴ-�i��,��}s�����@�oْ��Ȣ%VZ�GQX�W�LP�%}��rg�5 ���6�.��L���L-�Ee3�#��D�Ck����Pӕj�����W�+	��<n���s��u�Y2&�-�"pF9�����(u�����ځ,�mW{�3��M�*i�#V�L�� {M�8�L`l�ḩ���j�����<~��A�%U*s-r�	ـ��� ���-�f���D.�#DQ�u��eNCq&��k����Io�[�,@X�wOF��S�;�- 6P�{*�M�)A_&�uJ	8�k��� >h� ���*��B���(jE��Uji�'{�鯐���(+���R&��ƙ�u�#8.<��H�B�����Ә�3כv����F�g#�eԎ�ٹ�m�TRy�'��)��TN�Z%ߜJ6���&���;;&�����Spt�#�6b��<~�^�S����V�#�5Nj,E3`8[�x�3���/5	1[����T�1���<Ku?�3�r�G\��q�2J�[~�%6Rk�*�Yu��:��	F�i��?߳�H�� M�����HKH��m��ml�{:D�؃�����I�+��n-�kz����xm͸R��J�#��s0��T���2�;Z�1e���.�©�a5�r�ڶ=���:��Q��"D$fG*=��~���37����>��1�(�="Oٚ��F�Z�2U��=�5������"z��yl��b:�'Q�:̯�&lx��7�l����=�pF�z�k@�ӊ����A���7ҽ9[�,C	o�QyIX%�1�� ��4��1�x�#(�aDߡ�n�ช�� B*lC�br��|�>�Ц�^�1���s�
P�.�A��aX^�6�x�(�H�Q\?�����>�7��C\L���K׌;-.6���x��9DQtVW}��jq�᚜���El~[���J
�Avׯ2g���J�$����z�����Ş��[fX�ǲ2L�/U�޾38��}��"k~sȤ��;�F�ݑ��	��Z�x��s�xe'��{E��<#Wh�����rЕ�C�����S�A��׿�\���_�sT�W������#�"��P������d��7����b��g]����R�Q��j���)̌�Z�݃|npΟZ�B����J��yO�YՂ{��ءFW[it�������;�$�?�o1>"��H��L��,ѢC5�xR&$��ｘ�&N��������t�k�1Ԍv��Λ%̿5�'b-�ˣY����5��J������E�r����{.�h��U��6�a��0���XI���T��3�C���EM�7��/���$�2�U{Y���]��ejh�����ۈk���	0,B�}|6/s�5h#_Lcl=��n��w��M�
xt��
�Bk���9�#��+�a=�|� �$��l������
�KVЅvGe��^e\oZ���A<Z�q5u{۾�C25�
�S���m�- � <<�����p�s�ߎ�X��6As�_)��'k�c�H�[L��OEA�H�Р�8��`H�2U�ͱ��TąƁ���sl�d:<o�G�E���P6D��*[Z��O�aM\�Bw�%Iל',�_�kP��2jC	�֢Rg�*��+KK���wy���Y�����5fޅ���M��^'��rWIB]y�g��&	c#���@~R�(����B4-�{����a����ɇ1�Z��K��s�N2��Ar�P�f���(j����᾵�����!��ix���o^OΡ����CA� M����s�W��_���{t�>bF�ݶ��3��1\�6�E�V�y�����a��8;��V;I�y"�=�@�I��;��oW�m^�2��İ/�@8��N�g��,b ����W5�p;^����g�>�}��ʐ�4���ۏ�>�5.x&�e ST��mL;��v�Q�@�V������ �,%��S��Y�b00����]U'����G����-liC91a�Y�p��y��S�\)r����E�]}�]P��0���E��79�O�r�ʒF�/��Bt��Z�����\�{�
ь�[-�7,�~;�R�|���>=. _i(����;��r�n5ƅ�9�u�ʺ
'�܅�e�m�v�"y����`����u��V�*�o9d�z��� ��'Y���<��Q͠Y�?V���L�� ��n�wxc�� 'q���Z/l��5~Y��^[w5��ۜu\��i㵦�r�f�G�p+&���bt r�W��F�>�V��rp��'���_�9��a��7_��X���e颠�,�~n`�� e�@��_UMD��>sM�!�QX�s=�}��fpe%(�l�Hvxx��Q16	���Q�eQpܘ���� 0�/�80dWii�Ye�������A�%2�������i�Yʔ�c.��Q&+����5Y�.:�g�(��������1��^�=���e[[Y�D�=���������4��<O��,�)v��ы��Q����YZ��㲇{����C풇�³��O��j7�Z��C�+��Oq�
&Cp�pP�����d�D�x<���T�wRHU8b���(�K~c�^�^F�s��~�����g&�IO=�T>i�K/�!9`�eD5TR���;?�z��ǹ�;`2�D�|H�sXKx��\e��lt�n⺺�5�ϻ]	��O�3�.A_���O] G�/əI�m`���H2IaO	qV��à��N���Fr��X��}�+^*%�(3�u���K�g��Qk�b�Tu��������	�� 1��˖�9��o�(]��䄁zT�	s�LuI(�甎,��m�E�&� �����'p��#.p�$tl�n
��.�-ٍ	4��e,g��\�1�����<�z}6�?0�w9�}D8�ǑD�G
�V]��V��Vp);1���QKn>�."��rx+��U��R�Sv��4�z�2�Y�[�?%<�<E����x4�t�.1���c��p�]�WB�vȱ8�U��HJa|P�T�<�������]K$p�6A�#kD2S���D�Ҏ�!}���v��;8���R�'��^>t�o���Bҫ�����`F�~��-bD���si�D֪#Z"��$�r�{4��4�£��lu�����#vaN޸f���<���(��-�{$C�>0X��?B��n�����ߌ&i�CMIO�زYsASO�a
,ڨ�$���]��D�y�h�ox�B�{��%�)N8�r����0��>8��*�Sl��Z�4b�u��!ћF@����d ������G�K�cv�=�� �R������3�<HL;�dN�Dtd~-�I;ii��"`"��J�����k{r���\(3� `+��Dxg�w�́u ����!"��Q��2�2�9�1ހ����d�߄�h[��j�����^�s����
v��������W�[xb ��w�s��qnf�շ�t��|tK�����%� �R�$b�_����@%V�cA��������h�Len1:*��M�B�`|��裗��O:����I!��B|�e���~��aA>�DA0���y�9A�Dŧ��u@h�Ki�����Q���ݏ ����:�V/1�=�h�>������t��k��1�w;6$����nq@�s��4�A�hh�R����� ��n8g���֚�GB��H�w7�t3{�E$��_���=f�MO�7�F��z���;jnA�T�?�P(�����>�@yrJ&r�]e��V���D�Uڤ����'M��j: Ҋ��^& �
G	W�U��Ė�uF����"����<��#O\���;�IPe�rS��]�'Ę! �~������F��ôG
M�f_P
��-^���N��$�y�hsۢ~��R�kPE�;�-N<(0R�9k�J��d�T��˱hޛ:;cП?�S�$+���'W��8�[G�d�'C�^�+�� bj�	��;V���h�Q#�o����I)��F6P|��樴�R���dN+$bF[acp�z '��R6F����9}hsU���e�5U�t�Q�c��e�@1����f����0�Sq�E<.���<8}j�%������ ��q:8k"O[4�*P��Y%W������3CX�;����.D*��p!�L�A�QY�}�4z��G�)vie,�}l���vgQ	�h���T��{e�H�����:ro��`9[����5�	��d���i�w��A�!��Z4!��m,#� ǫ��Z0н�x�;5����U�3H^�|]ԛS��x�H���%+���a��`�,����7a����������c`��k.��Tj��f���*�[Q/#n&���������O���,�$�o~���#*���QN|��vtpR��3A�ԗ�nPE��*�p1nG\Uv����4���M�uĞXWB<��N_>��e �9qӹ����1r9�,��?�@fPw��h ��]��?˦5�����X�T�t�O�c�n��;9'̬T=�?A0�}�Km`��5|u��d�3��c��ԉ�C�diV��l2*��NH�n��دm�V��dU]��![=��k��~f�uK	���<�a����O�_�ˆt�3d�e[U^=.|?^Ʒ��{=�t�7��J\��Z�°��Ɛ���e����:�K�Q3�&10x^�im������ ��B9�E�2SWk��8��mb���,��3H���iٞ��s�k�6�.%jX��|+�FW��uuI���p���F�n�s�6`���h�ƈ�e�4�_��*����i���������H-��eJ;u��)�m��B�������sk���r�5�C��mE�M��� ��N.�g��W Ν�	�Hj�U����q�ƫ�ڜ�\���N�[c�̛��b&e�w��n���9�o׽�^r��Ӂ���UB����5 �.I��9_��R����闝�	H;*�7Q���IS�����81 ��oq��X��n}*oe�(��	�F�$*�Y�aJ�~�`�N%�砃|�l$�w|f��2�Yߣ�$��̿i���޽U����
��#��d|S����j%�@�Bϫ��r��x����$����F�u;��&;6��&b����l�c����x�9�l�x����򴛛��Aɰm��<H�rm+��<]�7���2e=�ހ���O�w<���]��1�B�b��~�T���i�z�*�)����+	f�s1���z�=��aA*8����N��PQ�/5�C����7j�X�Cr4�Ƚ��W���3������Ȇ����/��w0Xo�f��C�1|��H��=w9�̂�R�
'���Lڄ���Xo�����{��myd�/(�>�T��@����Ω�?Q�^�`U����^��xQ��V/��FF��t��<8���Љ`=Cc�V}��+���A`H`݌�c��=)&�����
8Ea�[�fOd�g��I����sH��7��ɿ�<�tӓ(���0H(/�.}Z�ݵ+�t	�a	ˏ���$([�K���jei��O�������o6�C�ZJ�e���q�\c��B�/����7�6��է��
`�IU�}�W}v��X����	�LZ<����H�܅�\lw�
�0����6�(�x�dÅ�dR�nɆ�7}����߽�d���0
�po�����*^�ٚt��{l��2����k�w�"���.�C�a2!�<}���6O({�h�ؐ��r%J�F�Kp?�����c�	�qp����AfS/��mJ#�V�	����G}45Ȱ� �BX��	�C��[;c�/v<V�4����q|M���^�dK�����D�|����d���C>$`��n��r�V՛�z�4\	;mS����\�
�=���Vb�C�T�Y�_�T�Y�>@��\W�]Px��5�v/��*�~i�'j{ﹻ[�^B�5��]�s!Q��]��O/qT�jjJ�*s� ��{#�â�)���a�D~C8p�v���g�BY���4`+�f�� �w�����1�U������Uqź�!&A����G&�ݻx''�P�,��?a�[g�A���N�<P��*�|Q���H�i1�V�h��R��TU���ړՙzsD�&�t�D�� ��d�쥈+sCI��כ��INM��IK�䶨��jwYLLf�Sd��(7,��p
O����Vj5:b]w3�⋇��gӨ��Aj�8��(��|�B�O�F��#�P�i�C� ¬��$���J�M����Ξ�����W���'z�O�bV�`���z�vi]=�ua��=��A2��m��&����Xe>�-��Z4��N��~�~�l�t�C��pY��p�.Ȼ�,�P�V�]��w//�"C�����]8���E����i+��\�b��k��7֟D{x�H* <�$T�ll�q�Q�@��ύ��o,�e��{�����\2�A�L�I�vҾ�������k�|B/C����0���(�]^��H��>A���j��E���T_||�j9�A6Uov�i��k='�;�x] *<Opw03�����4�-$����c�ۮ6�dGP	��;�I�3o(��j��d���bqJ%�CP��O'F}x[s��9j���B�D��T�1�&��F��v��og{z��|;G����Y���U�$Qi[�:�E�Kp��x`!q�"8�y;x�j�juUg�M"%Pt�������책MwNb2<EG�犋�e���ދF�T��(�SV\<�%A�S£x^3(!��/�od�@�}��g�_���6)ȶ���nV�W6�̐U=樼�P�R?�B�+ ��}I
i�����+�O�(E7�h�+;����N��N���%�����9EG���,J2�]� $���"���#�>���gm4lxČ�K�AEY�.�xB\�
��Ox���%�.��1e�����Z��u̶
���������Jn$�"[��;��r�3�����}1�v����b�Y*.o�`ۓt,�خ��ts�B�۶���`���L���c��XF@E�R
1bV�P�g�U�V^�����-�Z��=j$HEV�y���6�{f���pr��0G��@^��~���j��*�^HQ�M�G��b6Qt|zݺ��څ1ܪ�`֯��]z���('c^�W.?L9���-�GyU� 	R(M�s(�F����W�m�'k�wE�`�/G�Bg-��Q�1C%��݂�V��jQ�\1���k����伞9�@�J��ڢU�巅>��7�[��ќm�BfX��4��x��Υ���/P	�O4�}�k����>@)�����ITwRz�M��� W�~L�/ Uf�gȑ�&�0 ݛb4��4k'���uQ����{�?(e�,���Uh���#w��~����E	%j��)�f�g������	D�}y�mS�EUx�
�U�҃�{��|)&pѰ�� ��_־�Tk�5ڂ1����5L��D o��
����!�8R*EC]k?�b��i+�!'�s�0]�M@�wH�����;��,L�l�(Ҭ� X$߬!x�=�b��V�*����3BH�r��w��g��whzJ�h/��8[��WY�j�����a�&�o ���"�ح�ת(i�2�����hE��(~��,c�z.mK0�&sT__�2lq����������n���ɘC�	�1��<�H��L���-������XnA|��L��{��~A������%T�`���i�|ԟ�G�,���B56UW"����1S)NZ��u�AIyae�"Y_������/�����;&黼Ƿ.}7�-���;�?��6�X�~J���s�⼓ �!Q#��[��ة�e��k3��Oc�M�]��>�H�aՂ� K�P��0@��/G�R�������s�w�fݯ�P�W�j����t�H��i[#�	���X'�& ��7+��Q��i�!E\���ٚ�u��'QH+訉π�P�0�s��;R(�y�6.��X|!�`��Nz� 2�@���|ɀ?���0(1��.��*5!9Xa������E�|ek./A�F���j�mg[o[��T���E���Q�l0��ڹ:�R��d�?M�|k�:W��].�/,ΛR����H&���UTݩ�уR���w�����j}c�ˇ�	�/CkE&�0T��(=T�>�3�+�G#<��9͢��>%jcRqz�n��zm�n�v�����8���zf�F�g�$� ĜF��'!�QR��Km�AI�ޭ�ki�󑯗�Ь�����O�2>�W�gZ��%�n�Ȗ��]w���2H{``����.KG��AJ_��!�#�;y-O��ݿj ( ]��5�]�n���Ù�<�c�J�z�z\o�����ˉ�Ig���M=~Ff�C���C�#����%ۗo��V�x�,T�>�Y1�sM}�������*��Жa�X;ڈ`Q6�q��4��D�t�+{�|��#��c�8�K��X�Ŝޘ"7��E�{_����1���6��/�DSuosyǭ@Ej�����vǉ���*aJ�bh#�BC�Ce�-�)�Y<0(k�6�[�~sJ��tj\��B<n�V���L�����Xm�:;D�J�>Y��Y�� y�D�C3pvsCt���GR����J��x�C�-��ߣ������qo��[��S[�/m�dhw;4g�!�"�]Z�_�U&_��:�/8Zݾ��? ˼	j�
�󶲔�c6{_6LX^=�����a3�/�qlrJ�7E�3�O��f? ��$�@��=*$�Cw������ r+휕����DPP\lN�\�^���g���.z4�&�\��B=�����dF=�.��}�&��y=�����<�2ؗ��,�	 ��v�i�QWJXs�s�
is��-�/�\ؾ�=t��~S-�>��J8��F��bv1��Z�ꑜ.�߀�L�6(o/��R�b{�e��F��@����a�w������k��Fn�2?�9&@?�Q���=v^����o9�GBT��:ߺ���y� �&ٖ�j��b�V������@�۬Z�i~l�B��&me'�EL���b������W��yª��Z8��j�J*�g��ﱪ���c)�ڊ%�7I�3�;m��R�B�$��ֲ�3��b^!����s��g�s�;���� B(��Dڈ��T���|f���I�nVM��6�(��E�n���̄�i��(�Q>a�e>G�w+\�:)xJ�j�&�����o�_��5��ÖK��:�0o>`�S�5���	L�}�d��q�+ib���ӻ�+0��!Cً����,9^'[Wh�Qi�o�d2��r��@˼�1� ]Sq����v�ijG� ����a�/V��5M �5o�3��f{+�@+�������/�[s�j��r#���"Q�䲈tV�J�F����Q������E�܊Ɠ}"\�
H@{�Y�!�D�G��y�����yO�n�dg\~�c���z�{�������<JP��� U�E7�%�6�{
Bxz@�V�����I�q�w�ƸO���?�q��\
���ѕI�M4�������Fy,E�_/B�NR�v�J����zƓ�|.Ȧa�I��c}�Y�0%S[�P�ȯ�qj����?Q�y��C}>v��HD"l���1
��l�jԑ�L�mJj�~m[���K��*s3O��l�r��+O�S�ȹ e�y=\z���Qf͔�,@�]���/�Xe��i�/
��X�e7c+:)����Ѩ��c��IR�4v*SH� P8
�<8�c�ۣx�W�[�A�	�D���k�����ו��c��e�k#�۔<n�,��!&�����j�a��<>��h.b`�H�p2���Т�K��,��kW����y��ΕL=69\ļ���++A���<R��������?��rU���B�eh���A�$�7�C�����f:K���PS]Fބ_�7#3�j��� 4h�mY�S6��S����q�Ϧ����4sٴ�s�>+�@���5�q����#k���5%�mXv7r5�֖����<��LC�3wM�u�����P�ʊ	�y�~�F�o��d�� "�Au�z���#��bgI�z��%�X���8o#���ܥKu�1�_�H9_K��&�D&�#�搪/�]K��B�<��2v�?��(�	C#Ft:�9���J��@ �x�3��D$A��7�|v%��n���+%s ��+V,�Ur	���鹬��#�t��\����&��h+���e��gҖ[�2���.�"N�<�'s�[�Z�������n��V?���v�X����7v�ڮ�Sl��컅���Y]�h�8�����_��:�/�+2�P:f�K�D��@:�e�(�6{�]����2�[�dd�3���\����&/堝�?y�a��gT��UzOw�I�SL�IC��9�|�b��X�WB|��R��ˀ3^=,8�kb]{�%Zte�^kp̟����\n�(�������p`fo������vg0�+8A���f�]�0}�KrjON(��tvr�[
`�-��`3����T(�k��է��ئo�Ų��L��ά@��@ȱ�3]�ȶ/��K/,��Y��}\'�C� '3D��uR�U��O&sѧ�a(�Ƿx3�/&���Ϩ��)��B&�l�ŎSϺ�"����u� ��,��mݤ�I	��о��)uzF�4,d��$�hAbˮ�X�wA[�p��� q|���#鴌�Ž����44~aB�kH2�ČF�W��� Edx�N[��>�M/���`��`Ñ��w�cM��@�	sT�$��DEo:�L,��u?����� ٌG��]���~:σ�b�I��7o��:'0�uE��d�����}��gL]�v��WtV�C�5α�u�<`q�I ߧ�c��jɱ��$��gˋ�ƶ�����K�N'����_��<��	ңM1��*��	X��C�?!Gf��GÁ¤IA �\x�R���vH}}�������`�oZ&��}�!��U�E�F�#VC'E��Chr�+C�ѯs� �
�5/��m壨�ӏ�X��1BƁ�f�a =z^Im�USP��?@` 8�N1u&���(�k�S>aX�|2��㢜�ۨ"�~�f�%�`��~�]�7�3����r)���S:Kw㮝vp����Y�yII-�$\^�|�nT�}O��-��J��ZMڡ�AhH���Ҍ�o�-(,WY�#�����R�-��*<(jM��h���<~�<����0�6O�Ur֓�ѷ��A)��W4x�'��Vw�=zS%�\ٛI_�"mC�8a3����k�+;�세�.p�HCAM�6�?\���B��H(��-��KJ��ɸ0a���k�UMj��6|�3x	��o�0Ґ`k�b�%~�j
�������<�,~x��IB��/��כ�sAٲ�j`�d,�k"�	?	�=jl ��i�q���X%bDp&���o
0����}
?��F�����aU���7LR�q*.�˪T��{#��!���v�xAX0d�� ����HY��s����.c��ݦ�.�:��.>6��4�W{�o�	�̪��:7�m�Vk�c���Z�eSV�g�T��6 $b�m�Z]�HN��������7ߤ����4���:�t����Sk揬x;����qH� a�I���{����8M�-�O�:��7�[��|%�|B���V~�Z���V��EQz���V����l��m�|N���Q0�֏�p[��=4��Aڰ�ڗsj�ކ��hʜ}�ڙ�4�$���q`y�\��l���^2�vi�6a�m}O'e����š���W$��״!�,ua-���I_Smu��z,�u����3g8Qp�|�Ÿv^+��A�s1��ק*U�� �ש����D�zU������ ɋ��.Y{~�Bb�p:�P��n")-�_�l��Gv�fU��f��{}���y�~��}��}s���ٕ4���&L��pp��,����ϓ1f�Z���62�]�:�8I�!�ÿ�y��hJ������l}�$�8c-}N�s�@7	�皔�B�d��տ=髤9��b��_�`�Vd�J:�6�biU2�!�3�-*sDJ��K-�a�F���EK�r��i5Sf=����6�h�#t�\F����a^�mIR��N�k�g,��TdrX�����AQΗ^�ꕨ9��B�+mя�7@�!�qIG;G[o�����4�(�}jhd+^;�9��߅,��R�bSCX��7{�VK�����ܺh]d��;h�6[��CZ�t�'�@�zN.��3���ݠ�F6��I�o��o+`�hp��ƺ��^�Rp�E�gA�� d�x��vM�z�Gs�v����F�x_M M��"a�F͸wJ'"�=�4ڎ-�Y����5ŲGl�J�Ap˦\0/z����t�MO��Է��8��[P���<鈁�%��0�ˉ1n�ߑ�}o��� ��l�.@>2�U�e�L�?��0gJ5��x��I��<�2x)�e��uD���q���yU��9S��7�H9��"H���]Z����[��[$�l�� 9�=k�>W�/�å�RYQ�n"y���`'*n�� ��C���e����	@��	�co0!��I~<�̏����o�[�lXI�>�0�Wu2��͂?���,p����\�%j&0�G�e�c5vt�����F�G�������wV���
y�߆)�����<�GX�w<����G�RҖ�-��(��ey#I�#�g,����Ȩ.�«kDE�6�}���krs��sQ%>e�Č��77"5y��s�W]�(�%ʊC���ܣ�b��u!e�)��D�=���������I橹�[�W��좪粉?d.�V�Kl�F8�a)�~ڧƈ��,) E�o�-�ApT����n�l�.[Y\],z�㌕)>[�_�D)ڻ<U�y�R���DC�=�HK%IٿL��� ޷����>>)�k6"5C��+aj��P�5ȵ$5�X{'�,��F�V���I$�i݉�sh�|L��RD8"E���e���ũdf;�,��� �p����2�W@]�"ZD��W�dކ(���H��͗�Ή�oD�.yh,�``4	{'l`���.��}�OQ�ԇ����T )�,{c��P̐���9�剞=/ ��.��=��f�����4e�4�\X�\��%�����U�K�!��W鑹ij>Y�.�X"�I�=&�������˭�g�9P�.��,֬VZ�^at͏[G�؉#� ͅ�.�W���w7�v$H��;H2R'5t�$�[�V��|&\)l&ݏ�<�v�u���Z4a���� x�'D|���߷wRf~�{O�w���%l���'ڔ��T8���Жg�G|�;N�Qfv���K���Eea,!&f���l(�s��dHQ	�C;X�)<4��)��hK�|�Xt�8ɗ%l��q=~ ���jA8ćI6gw�P�-:��`��G�.���햚�U�uLVb<$b�t�[��2�-��� y>��*M��}�������� �Z�Z�SLk�*�֥�o���O'�i쾬�b���
�ٔ�f�l���)[�%!��W����Q�w�'�{�*�B�{x��dH<$��ŃG{�e��RqA��.��/�n�X�}�Oّ��j�/DmmU
JŪ6|Y?8�{��&y�.��t�`%eVO@=~Ո�Z]��1�'}#hB���Ia�C��)#K�_��=9R(0f��Y/V磻T���|�仾�=�ZUf~\���D^P���:�7�: �9���>^~��mu���O`^& 3�,w.}i6�;�Z�hBŇ�FS؀U������K e]��/��a���r��@�iՔ���=�xq��9t�7K��,o�01��6йн�ng�G��a��9sBҌ��F��m:��&&�/��v ������Z�̕V�c,���x��&x���P���	��b�v��e�ĝ��;�������"��YkB=���/��d�?��8��mc:�"R���d}���D���L�k�)J�H10z�RkW��-��A+�g���flK�F9�� t�&F�à���w���$M�"�� ���f��x�IN�d_ƌ�.n��WU�e��\0�>�br=�%�kUb4y��z���#U��r#�(*��/�/3�jxȋӥn�L��x���Ʒ�t�>B���P��wO��t�<�2�[XHRR�tȪ���Σ�W�p:�
uX�8�,�c��p@���?~. }\�ߏ��D����?(�o��:{�(�d��/,96�~ ~A�w��E�E�����>N<�U�����>��Tj�/<�~��	i֟֋�e�`�8����dSı�@���,sʂ%ʇ*hTH����jX}�%��f��M�MȻ�9�@��l�,�qm�CW�����.ᵄ`1�G~`q�x�ٽe
 �|<��X�H�j#�J��P��ȉ���>�<d�����ä"�TG�2���!��A�����D��x���ζ�}W�1p�ǲ�W4rd����!�ј����!�r�ޞ ���g�A@M�[;0�V5	I�ǼO�Od���|x��M��4�w���3݉�?bє�xR�o������VBF�<���F�}���/\�.�!��F��7k��z���U�\@�<G�Q3א,/�b�߀e`�v7&�����Z��!�/��h�G�^Tif:n�e"wG���!�s�k�?���wZY8�"��\ݝ�����O�H�}0Dl���@�7X�S}����C�@�ƅ�ד�T�y�MU���L\�\���╉l�`�C�� }�>��Q·�}�b�3M~�!yP���6fF�k�Y�hM�w^���p�}��<�l��oDZ��-�^�)\��zC��z��Y�&zxֳ<��y5caVu< �K�=h���Yxl��F����*od�x{�3�=�0�8�bz��AC!Bp�#V�ۥ�}?>���	�Q?���֭����5�����Q�FV�%D��F�'8o�ׇ��N�;*
����(+嘌�M`�l�口��S(����
�~�!�o�L$p"��mȔ�>z lS;�sK����< CAW��g{:ͤ�v]�֦I{$��Tmp�������'d4���{~{��~N��a66֔�T�d� |��ݙ�W�Mӫz*���.'ɱG�x�og2��Л�ҿ��׆���Q��ŗ����Zfdc�L�]s��V��[�X@bl����y┢�Dhus��Z����D�j�R?���.c���T�Q�YM��� �ϗr~�87Z���'�dg	�bH축1C6�I1ԛP�/pRN_�>I�̜��|$o����|�6ހ+���X��~���f����%2x��O.��20����"w G�ۚ�j�/�K:,��~�qXWֆ�I��>Sc@�şc��wǧ�;wf��t�6�
� M:u���s��'�Rܚ�G~��n��&l�� �ɡ���x��(9m6y'�ہd�����INV�[]M��=�^܏�)U�̕���֫��Qݕ�R��#X��)
����A����7�����}yu+�0�ܥ0��}�D�u�RX
/��e��q� �x�������epq�u�Om�+�o�[��!���3��x��qO1��!H�*v���s�4mH*Pu"(�۶�b~l�M�����d3�����_�,SJ�O�Q��2�D�_2۴Y|���q�%�y>�1i�q��_�x�F�$�T�tx>fwJv��9��#8מ�`�6���$��~�0`F�9�hU�"|��J,o�D�$�����!!6�	���BH�8�oV<��Xg|�3m���KE)��܊�<��:M�K�f���LZ�@�v�=��3���
�/�n�=޿�M�d5D&���'X\O��͕�9,�M����)ަb�b���mZ�U��J���\�������jh��;��c�lB"��S:s�$q��c�o`�h\���i~)Z	=�공�MF��$�i�O�2ߑ��r���]cE�Ӷ�Ebfu�}]�|���'�Hk�!����|�b�UӼ��'�$	�:-�4WJ��*nN��K�Q�Yhы�k��PU�A�������S;9>H$�_9KT
	����h��j�F�#���*����L��]-��ʸ����X�D�= �"rYrg�,:�^��(�̒�u��\Z��u���v�����gg0��גV�~�ıK��(���˽�T�?��eB�ʳ��|��2�3�US_7�d���$jd�bM�j�J�m��,�+��ۚ����ƿ-4�Z�E��6 W��1H.Ȏ�l�����xp������R�v�vH��'g�[�%���,���b���Dr�<���~0���������(P��Fizԯ|f�: �)v�p
T30T+S`��~��'�-v[�/���ՀLlW�'0�z1~���ayn]�)	���mA�	^k�����q	1�x���\?JpT+x(Z��L����x �A���h�f�5q�Y���/�r�1��&o��n���[���=9��ֆ/��}+�Ƣ���zk��d_Q����N������Z�	"��Ի�s]��N^$HX�`���c=⥛����de�a�tY������}��:v;=��>#+��E���u����78����n����W� �?�D��Ѐqq�&�I�?s'�7�S�}�&�/Ms��L6�e��}�"`���b��p����ݦ�˴�7�k���g�8�����6����x����ג�y;�$&���knc�]�Z� ��?�:��vu�b�n@W7�Vpۛ�c�c�ŭ������vL�)�Ԩ�'_�-'�������{%UpL��p�|*ɑDx�6��ѷ�@X7��`u���CE�!,�
���KR���BvJ��&�zG������Mt*��njK�4��(�e+D速^T����6ν�O�q��^֟M�o	��ǹ��غ
��]��6�����3��_5�1K����q�-��j�0��i��Pl̏���j������߫�Ԍk}J]mW0���h�#��)�.���\���58�CB���wL�
䋉��ܿ����Z��sh��@DEHU6�'5��1*�bcShO����G�>Y��J&g�CJVK��I��]v") vI����B��;��A�%�VX'mI�}M�%��B�C_��E�tf��� ��7���U%�N e�e�P��fc���[�y��1�dÌ�_���'��jW\��W]ߑ���i�_7q���~PT�b}�j������Tۤ��4������Y�Y
 ��ַ�Ga=keR���)dԦ���x����?jjVV�>*R�7���j4���>�b�ʞ�T��8���z2N�Y�q ���A��=^0��;P!��qݙ<?o�+�P��3�J��L1�l%8���dГ&�uqQ� B��\eH�b�N�^��gʚ~N�	�ا����c���V�Ϗ/!Һ���|~��jq@Z�c��>tx1�"�}�&d�ϖ2\K�1��F����^�>u�@�c#f�Fa�Hk����ƻ]�Wġn ���	�Q`�)L�CD�����?���j�P=��5Y[�ԳX����v=�e#�%	�RR��J��W�����V������i+�Qjiq۰$��[�<c�\\���G��R[��1ݦWJ�YL�H�l'ƶN�uڱI��u�D:����b�q��gL��Zx�s+��1��Ǉ��;�B���e �z�C�b^PO3|�	<zP�s �� �,3t������˻fI�) D�?�^=���R)F�i#8>�cE:MFJ�MC&���z=��}��"K�-Y�˱[��E
@oj㑢w5�ajA���k	�M�fɏmSI��v��y��[�������m�<��?�V�j
����������&ۤ,����w ��5�՟~�cz�y_�
V(F�{M��$,�x�&,��ᬧ�Υ�zhA������(��}�iq�M9.��Mw/��=����g�K��P�O�!u�E�]_��$Dy�u�!��E�A���X��t-ZA��@W�4��쾺�Z����7��ԛ%�w#vY:�[ܺ�[�d�۟B9|1|����iK�O�4Q	���
��'И�A#���y��L'�R�;��3.3�al/SW��T����8����B�u��?/1�5iʮ`&��n�$b! ��s��,����[�r��V\;l�:�7��:o�/��u���������klA�Ai|aY�!��-�xKs#o�Y��P�5�	h~�����q��RUFG�Ez����\�N^�S�&@��r�@QI�J�,R4����ސ0�=�5�N��9��Ż[�OI����e0NZ�#�������%_�X[w�u%�._�9���x�K�h�JLAZʇ�8��Όe4�}�r���ZGn���j�*9�.MU�~S����"$��3I*��xX5��ܭ1(q�_�/�,J�?� ��q�@�E�������z�x|p�P��`rF�Iź�O�QN����������&j���r�y�y"fx�E��ˌ$"�|y�[a��R|� X�gBR��`����2[o��L����Z��Y�P�@�]st=�B@g&Q
��{mߘ�)��B�u�O_��S������=�6����D��*r`f�Si�`���W����c!��7��FS/���'�-�����?����5��O�2�|� `��d~�A��EՁ���y .KP�=�"̣���'߫` ��2c2w��}p�dL*b\э�����yK����E�?z�� 1����2d6��\H���H�S��eMu�ӬQ��$�=-�yU�l�@i���*"A��-���!pH�hoܛ��(.�`r��q��?��3O�~�s�
X�0ƺ�^H�Ψ�y$Hb�(�O�)��s !r�G�7_��&O�8����^�p o�dY�M��l�!e��C>ug4-y	`.�!%�,�:��pY�^��f�
02����"���(E+Ǆ�X�@O�=��#�V�WӃ>�G��Xw���"tv3����+��9E�����!4����@J���\%*ޥ��L���Q8�8��>m/ڛGLȎ��H�(��,�5&����Q|���*B�Z��6AJr�j��Wh�-H��M���a��7C��$7�y�5QQ�/_*���
B��-)*Ɛ�
���u������;x�}����'�h�e��"�B�b��X�υTl]{��$d�����B0?p���tW���!Ɔ�����%x3|p�+H�K��0�d�cn��B�H���k�x�s<�e���O��_���A9�k'1P,�kן�]}�<v��MF�U�
J��z��g+�������V�h\���Vy��2�+?��Y%[��&7Btrm}`
�Qp�X��%�U\���-�@�"�#��
s�����=��	)wa�x���g]KCyMS�Lz����d��95B��	�FZ.QŸ 4��h�
'���2�ՂY��w3ȵ>�	�_ю�1���M����a��\�T��V�l�ޯĿ��#G��Yb�9���娄[��[}#J8��Q�;�)]��u��hq�tK  .�m��N����`3	f%��sX
������]���C}���=�f�d���{�ߕ	�ɵ�`��pS��}�O:	WA�����ֱ�oM+t��WUv�.�)�U�?lg�}~��,��z�3��S_������N_��v"��Ј+U�+�l�D��>)�&�Q�t�� �N觤}˨rQ|�����ݥ�;3:,�ʄ`x[�m�z�{���r׷��s��?ƙ��Y��,������;��s��1
��.����E[lr�?$�7�di��W���;u�m[�T� Bqϒ�64%9���?v��SN��]GI�f���4>�1P�fU��e��z�<��y��*�]������W\�ۼg?{64u�&��B�v��KRsfP3���w��kS��2�W�ކ�N�`(A�C������jJ9���U����Z,U������SvMA��:/v��єV ����/�u����M�c�5C��'�h(����U�M�zʚ��0��%�%���jv�>b�[���w
.�/���SL'��fA���)Ï[!.�[�L�4�-r�z�z\�O�K��3.z�=�D�
.�Z[���A�	�;lr�d.d�$���۴0@�Q��, x1��`����(��'4f�]L+�c��h�@+@��-n8V����=F���[�z�������a�؍�I;kB��ؔ���I^��w��}�"�6�lk�)���5**��d#��	�@��%)�f��8�<�����ϛ$��ʝ�� a���Q�$�nA2K������-O;=���w�tc@�A���u���3���m[�u�Y2eiJ��[�҇���d�/���ϡ8�����wY���yi�S��1�=
�3d¬�4�~�5�ٗ�r�x�9���;/u�3��&����D:�K�[j��	1_fo����Z�>r2Y|��u��ъ�V�O�M};¬��(�g��+l-�_;��β�#�s�8�� �R�@��B���L�Y����� 7�tc�=������'|�Pĵ3�{��*s]��R{��x�ո��yh����EFx��E-q>��&��._�p���xi���x���4)!�����<%'�5@y_P`6c$����?ZR�����Rx���>P����cQ�(-��<��<�X
Z�Һz�x�ɳF��8�b D�f��6���K��%�WuK���b6���K���V�MGP�ls^yRg0H��,;�u�������L{؋&�/
K����X����Q�)S֑  H������Q��"^hY�!vwD�C6A
�v~-�s7z��v#�1����M��)m��qݚd�!�a^�aޥ��9m��%��	X�8�vA���	�X��k^4�h���g�{G���u��^����Ƴtxi��?$��Q/����Ϭ��+E]�N�j�=�o�����-��9�=7�FhIq$`��a`5ɼ�[�M�yNe;H`��e��xX��9�'�Od�`���n�
~�<o���vx$�����-��q�ٖj=5�ԵZ6�-E:>��L�	$3���� �yks�!u��YA�Va���ob����5���X��b�H���~s�����1���k��X��J�����Ft���m�R|`u�����~z)�5 ����|���Y�=�̖��!c�b[����-\�s�ዦ�3Y��Rq�������0!R��FaI4Q,�t�a�k��f�g7�����R���X�k�7�Nj�e8��/�Zaǂ�J(e��M';��b��Qy՗i�yJ�j��V��kR��OS_�o��/���mz�����8��y+@���ה����~��P	Q�{�v���
H^��.��b�X���'�I|u��{�/9�h�]�%u��fA�JW�Q�ٸ8a�N{%�d������hgB6Qv�µ�M����0G��pNI�t�Y�S�yO8��*�s^����dn07zM�#�E+z�|( �xęK��D5}UF �f�� J��%�hS\❛+�q<L	U�ksͦ�36<��R'�4ģq�F�߾��[���\�=��<�9�>�Av#���[�$�E|���ivm�mq�h]�{�oa�ց>�NOO0c�U�@����-�z�i~�p���t(�)�7�5��s�(+	���T�ɀ�y`��0�a]���w�Z��ʕ��a+��O�0à��$�{� ���W����T�5������PŽB�q+{�ƒ���aAn�&����B|��4�QW������bL�wis,�	���λ7�7=�B,.C߯��� �a��B4���i�k���8l��Kɓ���u���y�����9�%��Q=����%A&>�bF=�x#>9�6�(ox���ce���76j�K[}P ��`6A&��I�	���=�(dSꂰ�F2a��z�n4�TZ��{��H�g���YF��A/ҽ�����x)�IB�(�
u�C�b<��A����m��7��Fޠ ڢ��6��o%����?7��
�AƑ`�?+�.�ZX8zXkg"�LrH�Zqd�u!v.�G7�H�T)����5���$��=���]�!Z�M$�
x��k�
�%Z�S~b��f�#��CME����7��+��j���Lк�[��0����JB�a
Աy-�6�*ֺ�߬��Rώ:�j��cV�S��	�5�Q���e����b��~�'w�jn�!����|Vm�}SEy������~U�(�Ӫu[�����U�Y��u�v
��\�j�����9�g�Uݲ;;�xߺ�h���1�7%�Ԩ��FVe���b��x~S[��3}q�;�*�N���7\Hd�R!�o��#7�p�차+�b{�SʍTA��T��R8s�$��x�T��J�K	Y%qM�8�|��j�M�|F�$�?uz��A���4�.�c3W䄢�#B�}xܻ@�z�'Z��hu�n�hCY�5y���J����.-�� f��3 Me!�>�W�n�3������r���$S�:F��r�����
�	��p���v~g�UFQC[D�aq^�u7���;<"۽�n�@)���[⃩[���hV!�D}����b���5�w����(g$f�%ZZ��:ϑS]������~�Zp�s���/�$��������Bj1�i\�� �������zp�8�=�=�|ј ��L�ß�g}�n���0�,�ö���qv6��!e��0��$9�+�veci�yB6[�Ό�R�N	���n
fC�YMfl�A#�ᵃ�vs��ba�d�����تf�6V��Z��e�m��&[���o�+b_�Sfk,|�G:��oߨ�U��:T��T��[�_�$�	gH��	1��B�r�6���O���D#~@��k�i�`��_&��u�~J�8����.WLњ��2�5�;�<�w����HPǡ{�me.k~g�4�m��{��$��%��u���Sk�/�>� N�����Eyd���uSs^��k���o�17�l%�q��Z��<��32R���!j��5D�}�l��ifi�D�'���P��?Κ�i�A���'s��tM�����o�V�9W�{��ٰӫ�ԋK�+[�yp�4�ԛrr8�ÌS���Zz�� �l/�v7���k��q��#w�J�S���E�Z�n�n���%`X�V�/���S_�fH�ޛ�rZ�>��hˋ�+D�D%{���j�1r�q黙�]rkG=u�5(����q��VV؎D����\�c��-��3��ȵv�d�/��.¾�+�+�~7V�DlY��f��훠V�(��6|����h1�&��!\�������*�� 5�c�@Mh��6Å��:�,�S��cj�mrɊl�ڞ��
��$Y�y���#,?AZB�á.V��x`�7�{T�cJ�,b��J*:�����F?�.`vKoxZ�~ڃ�iϢ+�x�&��Y���[��v���ڛ��]�0�x�ꐭ�E�z��嵃^���f�g_�±�S^�"��%>{��sW:{\��_|��Zȳ������0��Z>����'��)1wt�U֪e�����ݧ�����?[Y�h���s��䦾� 7|q,��\u'��Y7.O4�VS���r��վȓo��R^Ξx]�8�\�V��w�z��Ȓ�Q̗�)�I=��@���tV��]�*5��RՐ��A������44�f�G�{}��T q���Ne�>� 隗�P����E)j$MG?�To���?V���*��<��n�E����T9 qIw�8N>�[���Z#~~�l�4���	�4��>�O�%�����))@�B=�U@�oAm�ZL6[��j��b�O�0����:�NO����}��C�Bl;�ľ�ʓb �[���٣�l�D%m�������T����.���	�� DQy��vn��⼔�/�u�5�}d<�,�W`�Ai�thv�s.Q�?v,[f���8��bc6L;�=��׌ �Ȳ�ս��-r�0Nq�NG�D������m�-G����/P9V�s�_$����Pv�1x�)����R��?PM!�1�dj����,�p�<j�=Ś�i%@�X�4��	����F�i����c�c�sKb��m�CwxAeb���+�
�)6����<��8���	\�*�9o���U*�_X-r.+G�._�;"}�`��Iۉ	=-��9�ԻS(9ƃc��X����=�:=�qB�Pߺ\�M5��C��Ғ�)�C�os�m�t)���l��sr5�β#5z�1{�]K��-�}kv�h��W�}��e�"t��$v��ƱG^g�&H�$9} )��W�V�ƫl��1Q���u��on�)�����`�oI/7-"|����_U �[�3�6���K�/�g�Y1.���ʋ̟�&�C�������z�Y$��Tho�v���܄�8ڃ���iik�­u��dVs} x�� ��6�vO����U⧷0���h$�0!-��oM:6�j��@Լ��l�{�;Q���E�9V9!�^A�s��:��L�M��N>V��YS��]ȦC����FZ%��~.i���!t���Z>m��
ł	��j���B�
��=�1�{~���^3d)���*�	��|��3�^I�i�3�	�,rIҎ���y	#�Nʤ����;C��Gl|I�m����'��_�1����c��եz����P��S"���~�&5�c[�l���<S�RĞ;���>���J�ܧu���e"嗱�7!�`&}dA���a�l;��hz�B,C �6�Lr^||j��U/w�K�&�5(�D;5گzj$Īj�y����E#�k��GN��Ƽb��C�B
K�=&�B�m�AZ�8�_��:�!� ܉ o�]�-�4#@[-��!��!�)�ImO��qq���X����~��+)|�=�!���@��\����Y@Qy��%�R4��&lw�w���,/]묣�md�5�ۻZ�Mu�ծ������Ռ�&�+D6m{hU�YS�MR�3NO�mONe�*�uTF\�o��}���x��a���.I	o[ʉ�}kB��X���ًy��7�[��AY�D�:�d��,+}��c�=���� ,�����L���,ؾT�+�
n^i-�"��~�����,)����^�l�h��i+�җ�Or�_ �-�"��U��Zzhr��W��AF-�2r�%s }5S�����#0�tAV�B��-f�u���ƌ�sL�DK�4������@�n� ��yR�����a�(��/�4�1�p�8�eڞ�f>0f>5�{�V˓�>�ެa��I$1OO��*+�3Ȟ�\q�1М�����s]�k8��+�kSi�M��Jrg���m��/o �%ka�~�z�B��3pt�{��O�-y&XE,0����i;t�V�<l�h�%
� - ��l:�B&��M$���[�0���6�����TʳL-$��Q.G1��;9P(�ϐ��
&�č�բQ��������M%�]/3H��7�]J�ʥ�QbC�.�C7��\��� ƾ�ll=���W�Z�4)>O�3�PS<�1���xG�O�n���}W{qaq�����Q��?��uy���Cv�eH`���;�9Y(	#������ϘX�.HP�V�'0	�j+�ǲd.�7�r} ��u��6鲿���/�D"z�H�5?�J� �ڞ^	aC*�^O��=#;:ݾ��)pSNRcD�KTh��r;�{Q�I�x����[֤R~���WOu��UHţ���Fwht:m���DK����N;h�E����� ��q[�)�`�O�+NPL�_-a��%I%�!��VC��,G�m¢
�b��2M8�p41v��:���j�^t'Q�Wiw~^!�c�tO���j1;�5x��W�������&~P�\,�5�����~Hy���c��_�T�d�
E�{lX�@A�Y��cW4���z�L����Q��W���	>��	�2����u�\J�Lū�~�c�r���ׇ�I���
��G����h-ϕ#��8���H�]�"N�Q���۾�d�5%��)q�)��@�e�z*�G_t%�}���8T��G)�z�'תm���\Ц}Y�{@e'�!�&���I�1u/\>)�vU�vH y�+��Jf׿�׶� �M$�Ek]!B��?A�������e6O.a��ָ���3c1�����%��2%�r������H�����$]���Trt��IT(�r�/?Lf���c��5�&M{����]��� SY�b�o�**_-�g�Q�C��᲏
��DEhǄu��r(V�����]��'򤑤�n�h��Qԉ�)�n�潞�X�/E���y�Q� Jf��7s�)mi�Ӑ�1��P��d�Y�����^���N��1 �E�)���?� L;(��8VR�6~-/����q����&/�`��s�?��`��m	\�h��;f�Q�v���<��S�he
��Lb��.e������t�Ub\�!��xn|�I�-��ĕܶ|{�u4�(օ��Ց�W�M�c�Fj!����EM)}C}�0f�2����kt$�rx����mZ!���2�&�7f챺
N��s���k� \<툟�A�лa�|�7���s��J���$�-R�P�AFf��6Ӝa���̜Q,�Y�8���	�a��������F ��± ����bo����L���R��ކ����8��
��=��o@&+n��@kw06�=4�� Ip��H�݆�A>��t���%˅�22��k�o�(k-0�j�{��,�W:ܯm e������
���6厡��Xމ&o�c�����zwk��p�T�WL�[��d��+��d9����raR#A���G@@c�3�Ϡ���PlSr�/sʎ��~�?�W)�p&�s��PL����@��9���:d'Ye�Q�{�H�+�0��m"Q�*�t��x�M��Y�;+M��6;����P6�X��$���RM �ʚ�l�W�Ԍ�o(mrA顛m�L2q#�웽�se-��?��\t6�3�����gA2QR<I2=u�CVu�W�l
}Q����@�Zh�<��B���+!����� ;z�Q|'\l	1%��M�w�p��v�+�#����P����ʳI��s ��6�}�r�Wa��ʠ&�����5b;R��:�zV߅�8&#���mW'�(**k�(�3�>���6�Ώn� }L�(r\M�>�L����9Q�@J܊"����c	��\�Tu����1�S�"�)�)>����k����7��f)ZH�B��<WT!@�C��>�~'Ό�#Y��b���l +��~'�3���\�K�0��/� K����v���e|����Lf���va���i3��I�I�3�#�[?���� �S,N8���@���$HCCo�t�d�tS��E'�P�t���_.B�M-���=���ZA���dpQ^������j�X(~L���W4T��L������T�����q��,pg�����+��L1*#�5�i���Py�LbF��xQ�c�� ��� |�G����g��90�O���v��u5+n���o*/�Q`"r����sT:�d��y��d��&,����Ed^���Q����yQ�������:չD�;��c��A�}��ح/%1˥�@hHTy�A�n����n�K�n=�U���JB�eR�~ץ���B���(ucC#�Fm.P��斏[>\=$�|�=2#HM�F�<�+��ը(��>yJn�@3K#���^e�������d����k(�eNKw���m��\m{�����k���r��]�ۍ6d*��l0�Rc��JO���Y,��Lm4�#����� ��RS�e��,�FN���_pT�f��]���P��ɾr�l�}�x��j[�#��v�-�t�f���|xDd��>�2O����gv$4�5O��� �M���Ι��u�M��k�A�??�W\7ҧ�<
��L�����{A�:��G�"ؐ�����'���+y��.<�8p>V�{�@����g~D�-��0I+�v� �A�0�'�x)�4U��(^����E.�����I���c����#���]ͯ|�(v��P�Ӹ�10���H��W�{�|ˊ�BX�?�.�C����OB��gM��*��':̓��� ��,`���ϊ5�Z?~G��+`|�B��"��fá�bO�/p�sX���1��#
�8��&�I�y��kVbFK#

@�W@�����%����m3j�f�RZd��X��UL���SX_��)J	��r����xUP�ú����o_;QQ�¾�{)�$���h��	�`�Wa #X�Tr�����4�z�PX�YuB���%]ֳĔ:�ox�l5���~����^���=
��o���v��.4�p^!1X42���._K��~��ȖOp"xz��ͩ�J�,sjdq|*�n�o��\�xƤ��mҧ�/�ΰ�es��*���F+t�����M5Ӟ�Ik6�^�|��w��W�Ea���u��po7�ƺ�s,{�C2B�U�4bz��H��u��T�y���FgT�h���vҪTήJ3h��e���<v�\�{j��QR�b���䌑��o�Vҙ��UAZ�!�]4�!ހ�_�?�g�wa�"��q��s�r����/S���P<��P9� ߟ%Uʶ�<V�����w�J��c�2��␃=�a����<�5�$���v����Y+~���߾��+Y���Ę�Ό��؟��0�kj�&${�<��_\<�T���?�/���Ez�X�W0M�Y�Z}2���N�	��9쾊3����S�d`�P��Dy�IW��U�j�'IɃ�s�c�$�KY��E�V"�n&�woS�7Ő\��sTAR� �(�
��C�vȫjϋ�-K{�&I~q��s��WFvմ��ݮ������z�>P/^����!�!��te?'�	�h��D,,S�܊�{�)�6I1E���`�d69k5]�4idے?5~��r$�Ŏo��Rjwc�G��6=���V�����P~6BL�p>ˡo��L���]�q>�}n\C9Ov��(| ���j�
����|�Q���zF��$���B�Y,3�D�sd�m�N�p�y��x��?��:]��:��WG"��R|�N����}99�PY0c����a�������71���>Ӣ��Y8�T�
Rg�^,h��nv8��q�|�5�J���*Є���8�7�I��Oҹ[��_U�K�1��*(E�0X�-��LT�O�|E�����	q���|�(ѵ�Ծ��V�T�7�=����M��
aH�c��r4Ȑ�@�=���M�?0�u�G�K�R���[K����Ϣ�	/�6�~M)�W�Zk������B���@=�8@�o�&!a��Vާ�;�{�OlN��FTv`��}Gb7���>.��7Mm�uo�Ȯ^}��V�eQ����cQ��^z��6�@�QU�������jjֿ���*�JM��ͳ��m�T�@6$�t#@� ����]�`c`����SFx�,����ǆ%9؛���\��#�Gt��i� ���L�5�p[1��a�py�!k(�v��(��B�̋>�$hXJwL���e܈pG�ִ��kޅa׳7n�x슛>�%��\��$ Iލ�����m	vf�r�oN��3�����k�����΁����1��YI�A gXq�9?˽9Ul[?g�bBWS��O��v3¥ءӥ�{�����dw��&�i���w�G$�w�]����g�yտ$�AmG��3����S����|��Yh)rn���Ept ��?
z ޘ�
��J��o��+�ϻL�r�	d$V���!(\V#pe;L_���eڑ7r/����샰�mr���� ���O�Rh��`�QZ��1=Y���F������L�w@	H<�G��W+#�x N�4BA���{���4��OX�;5"�]��M�wM)�7��w}q/ 9��:�u��g@[,w� �O���P��$.	E&����+�
�1ǻn��{9)��$Zg*��x9;X�����X���=��i�OC��*��h�~a9���'"�U+vJ�,��t���\��n��'Fw f"�Fʯ"�Ks�2��I��N���x#��1y7�E`|긻ƿ9�r<��8y*x�[v����?R��dH3ϲ�c���I�����mX9��U�v_V�Of&�}���9�x�WϱBt��j�\�y���ۑ���G���2�י�>#n]�|W��f�˸Q��pq
��#�ݜ�#�l��O�Wh��7<�ї�>�bC�Ǐ*�a=}����^\a��!�Q:�Ϳߥޗ�bF\��,�8�@͆��vńۗ���+\|���A�Ʃ�n�6��Y�����יf)��������[��,ٔ{@Ϣt�B>QˤeJ"pO�����Q;`�F�T�7��訢	��j"��]�wҏz�k�Z��q��4?XI�fM��uAW6�I?�1�5�̧���9����cu���:ꖧ�� |�Y�_%xW�)u�vEϩ�g�Cä��#P7ʳ�k�ܹ�BU��kt��-@�Q]�{ߥ�
����q�}r8N�T�^���i5:�tZ�C�o��U�����ጄ�^�|���+7r���X�=l{E�tz(@�g]�~�E�l�h��E	��.��Q� �(�n��Cb�T:^���=����o����N��N�_�JP�#b��݇5�8�-/�S�}��4~����a��ۛJ}���[�q���}��}�v���x���*���� �5&���zG��R��d�zmb^L��Ǌ��]b�D���
����?�(�x�^��}��N���o����`��D?}�3�_p9_�9	ք3��!�Y�n�8�����T�����|�v�S������5��E��!�Lo�E�T3D�{9\��I�Ъ�X��a2��/���;�K�C���ގҵ���-��L��Ҹ���^Ev,a�������3��w�h���."�9���+�j��7�wO	�N�����,��p郅��V#L@8�BﱸOn�C��׆��p��-H.�L���&�pc��G1���n�:"��X�wEH�׭<U)�z�<�f�I,v]}�ڡAV)��8EY �D$a+��	�����gn��Y��t&��Mf���؇��R�
���T,���t�*�;����VI�65����. �g���9	~���n$ܭ(cj��`�P�LP���{�q� ���x���ƥzB܌��@u�c�Y5V��p�G(���?�n*�/�x�E�b��<D�b9��]���3XQQ���6fqU�����{e��H��ķ��5���b�+9��Op��9#"�wE�!����*�է��L�*x��R��Ȳg��&�3��k��WhQ�C�!�Ґ��J��^��<��C��߶��wV:M�� -W�a�y��t0柃5W���F���l�[N��f�>r0kݹ�	���]�jГ<=��MH�m����kG"k��3�k����m�����K��渿;�mvIȓ��mӂ����9E�sky�`b>�ܫ�qvz�FE`Q�W!��C'$wY�$����g?]�u�:"�G\�	ʴCB5GW<��;�Y��Y�0��,���q�xꨬ�S�!f��)h�g���0�7�g+��M�����������Z�ڴ1�U%������5�$^R�d
N��i�y��ֿ�V��|c�r:M��a�N����Sv��鵩�R� %����&�Y?n��S7ΡnnR"ڣ��E�{��e"�׋P�+e�)t��Sq*j�=���?�) ��I�D��J��ܟ�5%����'�T2%f�K 3��0Pn��y8Ό��ӛD�A���KU/��uk�B�Z�??>�%���(h�q��J�w�w���`��ݞ�8r��p5Y�~&epГ>w�*��e6�4��[z"���B|l��EZ�ӼX&ѥ��k�h:�N.&�s�|��PL�[��_�{����������7s\Vᾎ�bi�:<-P�1�fc�����*j6��=���Ӧ�Y>H+}��~1�Fx����󅦋<�L���m" ���C�i�6�t5*��i� _Pϯ)�N�l@���иf�)|HO�/%���Y)��d=+��٢�α��|�����뉽���`!�o�)L�d��-H�l+3��{zq�����.Z̊n{����:,��'�}����7h~}q�n�[RN�l� q�x�ȗ�u0�;��N׫�7��e��?3�H��`C�>�}8�#s�؍���>�l��-Q�x����D���C��Y��Ҡ^�b�]�N�Kp�ή�,����M�膣������/A��){�R�����=���%��~���p�y'[];�6���\�mH߇t�	�+�t��o��A��ae�� ����zn���(��������Y��(>l=�S̶֝n�7u��-/��Ӆwb�ŴP��������o�U'�`]ɯy)�o�����U_�2ъ�^�Z����hq�>�Ns����\~$�?�N�������� d�7>�8N�Qbu��}��aG�U�x�i����,�ӝ���e�y�]����d]��t��9�� �"���R��s�o��R��@ݞ)��^4�SY5�Ҧ��S����h&�� x����ޅ?b'U@�$�{Ӣ���Z���w1��@u����}|Wd������ă?|�7`sJk�Ԡ�O�����H�*7���Y�\�C���x_~����&ɚ;��I�����"A
9�EĻ$`��<V���p�~�d�.>�T��d�	��_���Y�O:�gD���@�t,�m�26Ww%�\*f ��p|҇*Dw�Q>�������<��ה���6�,Ptb��!:p�VD���AY�����S���xB8ֆ�.�, �����e����4=u�j�K*�@4ص:��*�$��}�A����\����v/�"_R*�4\��X�}��߀�H��e��)�BÛ/jh��������ZL�������y����&&�æ���P��X�V#�Y�����迊֍1�VGU����ίya�? �~�oA�S,M�"+����4���I#k�}��I\ [��~�0û�l�^a�Qz�X+�2��{Es$Zh)�a�F2�¹�˨S�nhǣ}���� eyv�:?%0�E��:�;���GErXz�s����,�&����~�� N��#ayM�&�q�V�P�]��Z�OEuKQ�0���̖$������g(�����E��~ ����Vn2Ϻ�Kl�7�jG��tm���tNz'�s�d/�4B #G��Oh���6�:w�u�����mq{T�_L��
p�R.~>�I��W�@��pW��%ɶx��-�F[�.��#��yFƇ��" ��B>8L����ǵ���Ѳ��70�"�Ѐb�%��#���$L*!-�8���u ho�K����p�&�#��$2�%0�G4�Ӄ}���Y���HoA1Ҡk��އn8�W��JH] {������)AHRc�k���#�j��'v~��=�cB=�b��^�Hq��ҕn�M�sl���g�&�h3�A*XD0�N&�hD��lz���v��&�ƪ̚��m����sq����=����y �Z��y
���"�$ۃP�|��;��+N��^�S��pi�/y.�]}����=S�J+�C�� Mȑ�˴�t.8�d��	c���ԡ�01Z�3���,{�%�=J�$��m��kSj�9��(�J*�G���l#��Y}aq`� ,ji���7*�#d����:=���|�[����h���q�C���k�?/궎d�L�=��q�!krX�4we�F4�3�������Յ)/Ć��`��y��=�P5� 3*��*^�}-W�	�;^�ܕד�|u�_��Ǻ���@%�a�$�(u����c�n,$����c7�[���x^����njq7iIג!��S��5�By\]��ϵ��-���iB��H'����$Y�;��XN��l[�Cc��>Ms��Ŝ�;��˪�1����N�R^�Ǔe�5�Cz�Um���O��d�_��hҲY��/�Bߟ�^����Z"���
c�ᰛ�[�s��.a+�Ϸg���w�8����(��Z���#��4�m�xC(��fi�?�HХ�f0s��]Ō��Ʃ���Dj���o3ܘ/�.YR.�ζI�b���ƣ>=z�-`Mu�,�9�N�y^�$�v�k���<t�z�HzF^yv��=�( ��Hd����p|F&2V�U/؂���(��:N�a(v�5��RԠ���׺W{��B���a�r�2=�5_��&k9�c��)����������m-1�Ð��> ��� ��g�����0���B�\h��{P��6�+���Ȉ�64���E�-FF16�Q��M�ې6m�YV2D��\�Z�{��+��bMe�>J�<�����1��t���ʻ?)+R���6E���MK�E�z�r�'/���kҌ����Ia��L��R�/m��nn>`�i����!`�"K9���	�OL[s�[�ي#�6:M����/ވ�q��Bͩ]��C�U&s� ƑMrk���tJ�f�@���/gH�B��6�ȏh��d�N�:wI�u8,ݻ\��k?���X����_�b����e$�R��ʵ��5��(�EDZ�d�868��]J�hp,P�W����V�ʡ���~`y�p�
�t��D>�,�ڋ��/l��P	�L���s�zH�x.��>II�/HJ@��3M�i�d�]D�<��WV�@�i$N���M���Z�Y��s�i�.�������B��gʚ��J���aI?�����ֳxt�uC:H�K~S����յm�hM�G�@��JeQ���&*j�_Ax���-�#<'��k�;�JBvl��A�8h�e�2)�v�J7!��3��3Z���6"�I�A�b=@u�)��e7z	�$�AI�l�i���@-��8�@z��Vտg�a��]��T[�3Z'�yH��I��{q9Rm���C��\\uM�RK�5�{k�F\�|.�K}%Ȁ���!������$�I^Ur��?m�����<��wE)js������D�VA~��t O��q�Ln�@�O.;?YB��~B�a�� �g➸�n�2DwV.� GPY���w�Up�M�8XIS���H�c�'�6~!Į�`s���C$N�\�����������T�l9rK�;ˣ�V�ީ���,�
oW8��Ҡ^ԗ'q�#��:�	�K���Jśc`��
��~�S�fP��)-d5�"�㦔Ы���C(�N��8��rgv�
�]�C��r^s��;d�.1^�Q'G�?�>�^�I��6�T��5"bc���<�N��Jm		�?�c�P�r�:���~�u=1�5����`��]R�P�#䣵�� �QT {*<�B/�uT��>,o�6�DW=b?'QЦ}���w <�W�8�N��{
��¦Z� %:6�����d��L���h��:�!N��1��o������OBB��Ʃ�D]�|��&d��nF����I��+
���exL�����쟊��oRk�-ħ�
h�������(�ن�����]W;R�	޾h;݃�6�ck^M*��Ֆ��67KX�K3����ڞ�l�~�iR� >�<x����D� ���}����7��N����qN?��悈�1�']B�s2x�Ќ��.?"�a*2�~W�Q;p0HG�}~�yx�<������aQ���L8F���W�����vRu]��9uTu޽�|O��@pb��)P�O��P5o:�v����2Y9¨H@�*|I�%yPA���4e�=ȳ��6{���dC�%�:�Kizߌ+�Um�I�^�jpT��W�����x6̗N�|<��ʭJm��g�{Si/�N�C�?��+|��烪I4{�Wx><t��"��gGV�?oKy�+&�kB�p�v߭�!E�f[������U�Z�6��#�ηQBFX�������Ђ\X",&0L8O2�fY���<v~�b��{ ���C���iOl?��3��6
����NuV�X�5���W�h{0���6�g�Ԥ�x���Һ��G�so�,�W����Z�x�D�B#����(��Dk��������$�=�����C/{�S�#\���ND�j*2Y�ѧPR��z
�t~^_���1�A�	<�9N�� ��e�t"޺M;���f�fS�e����Ȏ�W�_�s����wlh27A]L�k.f��(�6�h�a݀VQ$}Lg?`g�$=%� ����4�O����-z�3��_�{���0Z�#��T�@��x��޾��T����XM*L(�������t���rW��s�>L�B���6m���wK�ų����V��`S�1��(c�Z_�C^��:	7�G+�p���j�s�w
�R��"���N����:a-M˶t�DM$9�����ߓ���kxr�֟2��2�j�
�������L,"]1P�,�//_۷��8�4`<xN�[5R�&n�N�PPOHI�,�!K�i�j�*���H3ԶA���O`d�0q�����P:����O�h�F)�gM�'P(���i�!�P�+Ɂ��	O���Xřf�&l�)
׮�8	`���P�u)��.�i��pԗҋ���|��2?��8����B\�<� ��]��m�&��h d�Vd#{��L��y�/1��J��@8���Tl�|)�w�X�� iJd�f=�9��v��gݺ��w�=�Kc ��D��g/Z��X�$@�����s�`V�g~1/s�d"f5��AH�FNϝ��M���,Z��Ӆ~�Q����0LU|؞-�'ڤ`�@�ꏵ+�W-0�m��0��XKv�}��\�U���չ���!jSyƳ}/�s�Q��ˠ�dj5�d=�u�O�DI�i$���	��=�%�(FO�&h��z#Փ�2�^���%���i���D�kOw����Y������`2��r"��T7i�,�K<��66�a| �ա?�N���Z�������E�+֓���bZ������U��z�UJ!��CA4^ነ�:�'(xJ�7�~)�aαZ�Y��+����ո���68jSt��j���G�i�tW:Б��UtN�G7{[�<X��r��A2��|_	��wכ���Fcc�_�(��V�������b�v�Ӫ􈶨?xՉ��C�}H�30K�!P岯��ӷF?�ۅ���"S��k{s�0�Jp�xM����Lu�ã�a�@	����g����� ��]�f�6Q}}IU�7�}_��혛%�3�vH1�@�`[_�<tK�(E�8܄��%��7q4̴?F�E�lu���p� �ǻb�����;��G��]j��הxz�'J�WK�LЗ�)��q�*)��,6{;O72|Y(C΍g^�_��ZsW��ԼN��ͷr�2�O�Qe?�l�eD]���ȽR����
v⣍��er�صa�fw0Y�x��+g�0��A��a��n���q���w������F<s�;�;��Qݹ�TK��T�yMo�"��3,��<E߭.	;�@��i�Πo�2�e�ɻ��;P�(cF1�Uƞu��):��~ρ1�B���M�{Vw�p���%��vb��՜�F_`����[�S_��~�G�,$Q���fn�F����5�	 ��4
|'@I�%T�.��}B�鿚y�]����c%6��V��R˾ͅ
p����L�� �bܬ��[��n[Y�܉a�@��q�ނ�sn�ԓ����
&����W{��_3��`�/3���f��۠�%��E`7��������L�!W>��5��6�dbxF�W8�� 6��%���>r)��T������(����u2]�n2Mj𦒗�����*�o�N�!��̺I~���(���}���)�<ȅ���J��\;�{.�/�a$�ϝ]{I*~z�B�y�Ƿ�Mo?�;Č2��GYkP�鹻f$�� �)���P��!	�'���� �>aW/+1{3[��E�g�%��9���1q��|��,�:;��Ig!�p�R�ٟLZ��|ٮ�%u�͈�s�w�&�y.S���<H���;1�CG���c+'t[�� WO����;Bx�>aq|;�An��2j��F-jBz�b�����um� 8gׄ�D�+�"!>�z�������Xi��ת]�|��m��Wt�y�h-ݽ
����9���׫ƛ���J �l5�$m3�|��A�q5!�O� � ��5vF#.������O�:�BѶZ��h;+����<Hj+�2ɂj���?�ʄ �'������d�8j����Fʌ#�_�YU�f�,��o�Sv�Юș��mT�l�2.�X�]]mB�����4X��<�J��P4���<w?�����ڜ|�W�~�ejVڧ�<"��Dŷ��k|~}���c�p�TR��mj�Ss" �D�D8�SlzB�h�ن����$�u$���J|k���V�;{$�*������K��z`�CD��ɝ�X����+�,I1�*�hd�R7��k� ��DX6�֗�y��C������>��\�b+$�NB|�x���-u��v��@�t�����a���	������ټ��ĩz[��؈���,��L��zw$�OV��5§�}Č�V�<2���dG����W�l���
	{��S=�rpX|$�w
Zõ-gz�N��ni��[5o}���2����^aOj��'x����6���>��m�1Ť��A�������0��F�{�7k�<�N�F�B�Wq�[	�*ȯ�T&�jX�Dʋy���7�x.7�ح&:�|���,������"!�sYR&1A�F�P���h��i�z�Am���~m�B��'P�$�k���ĎK��k��⏆���![Z��?qL�2��J|����$��TvQe�B
�V�vX�R�UJϫ8"�#4�P�UX�j3x��}�l�A	�@���H�)&���Rg�'ڌBl���+��WW�%�,�e�`������p� �qL����a�9�dn��J<�;�'��K�wE����O����~�[N���W�<�#�����K��O��w�V@�����L�_���^-*�������s��:�#6�1О�&n`\he�������e|��̗�5a��8���r��=��T��\m�c��"�#�� =L�lq��/9�� ��~eï��,_���|�A��z��dX�H�~oL�JO	P��`c��j�9�K�߁��ǹ���簨��T�6S��r��x_�5	D��U�1�{�� y�LM��-��p���;�i1��AyL�u��	!�]��������H(��S�R�J�\U6���P����BeU�²���=��e��$p��(�|��ԉ*��qj��QʮٝL]p�岉�^M�U��|5L%���CM�y�{:Dˡ}|c+{z�u�=������ab������~E��8ĴFՌ��L��m�A9Cڊ��zG�I�q^���0�	e8�����13"h����T�WШ,�}����(�t��{��]�����F��u��gS�$L��C�'>H���b����x�>ˏ�����C�l��m�˵�gp��wȡ��֍��Fy�C�Γ!Es�M[��ni"hM�eKK��8J�&\��&����M����/�+d��3�Σn�xR|��I�.��j-�mp��F\զ�9tw��F���ޕJ���Z��D�O�(N��z��<�9�]����W{B��������o0YkxEP�'�<#�Ga�%Q��9N�w��oYF#NJ\7���:+:y�u6���W�-�}�A,KI���:0K�ߵE��h��Hv�!�1vL���o�3Kk�KE񔼚#$��cy��>��I���x����-ʠ�IǶ��sG�_א�)����-;loG�]��t�,[5�G�ʪ�<�_�`e�`�F���y��3�2�����P�l�;����~��eʁ*[7��S�NB6��������}3<4�ﻭ��<�+�W�k�&��*u�jo���ݨ�b��#���#\kmP�=�D��ȶFX���`_�O���Fa�Eְ�8n�s�B�.�7L�q�8.���w���m��{U��@�z���\��$I�")c�.7%s�.s�b늯h�, ��D�*�Y�pfl���Y��]GJ{Aq��MJ�����77-l��|]�'AS�N~���]ï*J_�R��=5�\8�"xɉ�IXquLOK���M�*6\�#D��r/]m�*}� ��U�bv�r��ɴ�b��
R�݋�ȯ%�m�Z�5��:��^?�<�wl���o�#�{�Nw�2��u�	~B%���4���؄�V�#�rQ�>�,q�8(�����EoWw�^��(��CҼߊ���
=S	�`+�u ��'Z�;��� �P����#M��D�e�
�;!��/	�W���%���c�Ž��U�N %L�1�p�CSi�ɑ�2�H�NѾ��g���aPo>�;K��*��Α?5�9%Y����|�7n\���A�s�ygr<+r��N9��!�l�󃭟K]
�wT��v1� X��,�D5?L�N�#ԍ�� ��!�\�n+��,�JC��ã;�6�#�uD�c@TXY���F��m�,D'$�r�\���a+��W[�s��$��_���!c�3���Ѣ*�*1�ܤt!0�%�H����mI�L������<���ا�/��5�"]�Ӿ�DȏY4=���kf��g�&� ����}M�*H_q;^^��4u����LY��N`S0=�G��:P�wYA�e5�ˡ(%���J�{ҡgnM߹٘iD�@�L����?�f������v�S4�*��(��9��n�AMd���F.!S��1t��F6��}�.ZE�\Z�����|���y`L��#�`��,2��gD���������3�cA-tN��rs�1@�E7ιT�[�I����!�H�߮��{� J?Q�ܗ��,u�d�_U�r���N^��9���b��T�&�Q!�H�ũl����1�L��bᕞ���.�')T�s�k됵� �yu}|�a�tFK��&�h������8��������o��T�Mv�n�)˽٥_�F`R�=H��;aG�`
�/��K.�M�\�m���b�$�2� Sf�\!⹅~Z���Sa���HFhO $��k� �g(�R���y���e}E��Ј3�KA�\�C\���b�/�&�ws�;��ز����G]�l>�Y۪+��c����7�����ٽ�8�z�5%�v�v�&����znY�0/���u+Z@��c�1钀\k/��O	�BZ�?�P#�����"+i�x��a�s�c�G>byi�)˭�%Y ���}��,鱮#�e�0�M>�D����_�D��׺�-R�.F@I�?ھ�
�u�Ϊ"rk�Ǒ���-8T+��ʏ,��9��zt�6��Q�]�p�Y���aZ���yu��ڑ�a�M�O����KY�/�J�W�=���Q�+��]3�'��ZY�z��ݹ�ɉ:G|��ҊӆNa[B\��Iq�/hCY���S^}O�U�������C�>*�O[7"�=o�pI��K��E�����ޛlM�L�w����=iI�E�r��<�J�}�^���ye8Ǔ�O�`vS��%g_�Sb�Ql~�:x7��$�����2���]�q�����tH�Nc� ,������������c��+�pS���]�I�M�K3�	��R�K���P��[s��fX#��f\/���F�2/��6�z���Ĩ/9j)p-(q�����)d�-�vq�@�r�%�@�.��R»�J�(gh[�1H�Uc����l8	D��Ѷip4�����ӂ\:<̄;Ը��gj��SѪ�\��GI�G���y����#��ݍ�5I�[�G���,���[�b P�Z��E.�YO0���/�O�V��UL����ӯ���^Rf�:X������)*1��h�-,Jo=Y�H��;�˙�U����īx�Z��ˆZ��2��S(iЈ�BF�K�t��9�/��Y�$�,���R:�͔��J��}��qr�gz��VAB�8o�t�b��!����BI�\��r����ڄ�B\�w���e�W�1�c!��	d8
�W�GFSdxӴB�c+@�4�f����bxwz��Sq�PX-�;���)��٭ˏ �m��g#�����5=�	���EI0�Z�Z�9�Ү�G�ϲJ\I������`.z���@	�qt�?���2��1YW�qDa��"��T���Ψ ����lo�S���M��6*a6�@���g]^�bAF������o׵[����>�!��2& �4Q�Ae�V1�^L�(����
 �OK�A#�ŊG�8����]Qf��#�4�h^r7�D(�/Kﺛ�E�]�Fe�7ZfM��"LG��|ނʺ�-O$��l��l8L�QҦӻ�<�[�\�~7�=!��N�^�4��������[q����#�($�Ra�:|���DX��׉l��*�w`?wB~�����^�	�z�9%V�R����A�S�,u���P�tK��^}�g����LU$�/>d�l��iT"�q?�>(O��E��y~p�-��e� �{�h�n2G( ��	����E�`X��/�!Q8��q���`l�Gޯّ����7{�^ ��l�S8�"��"��'g��hO�7w#:��9�U���(�f�A�n9�J����C�RV�)[q�L�bEi|b' Er/��KW��Yց�)���A%n�2�8��y�v.�.q�@G����Kt�f"�2���G���ɕ;!^��e��C��+�.rwʬx�(�{�����Y{�����������6.P��N��j�D�^��~L������*s��� ��pgu�ؕ��x�x�;Ѭ�2�����S	O0�yWf�Éۙ�������������V��j�)��S"��y���+(!qD����l��j
y�bڣ���N��T���܌�/�-��~A�[:;@8I�>�Q��ÇN9�33]�0�,ȍs /�Y�3�b0`�"���V%#��������D�Śh�=�ywȸ�|����K%Z���X����'n6��I�%&F��'3
i1�H��m�ߍ�&���b�^)8.�����������9�E���Ѓ��V��;�c�`����j��Pp��o�=��=���so͛Q��|*��x�!�T��v��N�M��b�{W�f�]�W����Σ�L-�a�����y��{�]+y���:�7�=���)��3{�ll�lڷ"���tQ��np��NjL�L*����k]�,��C��D�����&�~�%f�`j6��I�墡t�إ[���!�kXv6���S/�P�:ԊS�}�x��,v8�.��C'��?�Pޕ:��_ī����tq���j3*��F��J
"R�_}-,���M���(���f��`oK�Φ5d	��F܇���T�c�v�ҷ٠��������X�q���lV�U���X뢗�^�w)���U� 5P>�vqLR�:�����;�Lѽ?�Jfb�j��gHPlA��W�\��V@���X3A�|� !��,c��"��F��l���y1�Aaùd���cf�whsut��:IsLx�0���,��t仯V(�5i�i�o��c��S#���G��m�mE�DR#�V�zEF�X��	i1��kr�K{���bqꏪq#5�<"�9������V�r���_���z���hӣur�.ǕΈ�yr����(J�o,���x&D�I��{;'߂'�;ejx�E�2�t;�����L�'ʞDJO3+��E��xϜ�ELa��a-_6�Ӡm�M#��vS5�TF)���R�wh�B°��m��Y^̱�v:��4��6�o����(�1 i�p�E�+�_55�6.����g7Jܯ����@��U|ʙڹZ��L�?�<lg�)o��<�,j��Gl���m�)�PYxx ���w=��͎[E�h�4��`�����r]9ٚ&�C�e<�c��w�W#gb�r���CV�|�������؈�UΦl�h�J�{�(���T}>�ש���h���cO�P'[�;TMX̔hMI_-������>.�KO�
���K�kY��l�ݒ�ZǗ2�W�1��ּQ�{��.|��wQN
0�'�:�C�!R���6 эX���!�J�/w��b�-ч�f����~S66Ѩ=c�	���K�{�,��Z���ѻ1��U��1ݵ��@�j��\y3K�� ��{V�?�k���(e{��h��jKQ�#B�-�ܹ��T�k=���Z�����2��fU�SP�d:��d?(��L���Գ��7�vq.i�Oo���)����Ͽ���䚲]ǰ���0Í�N
g�DJ��SJ4�s_�H��D�m(�CuGp�S18���X���c�&��][�QI�����ޙ�<l�k�S7����Ծ�q
��W&��vtL6��<�7�R�ޑ��ݙ�����K�sx /2WT�|1��1��lA����#�5�K��{�i�]���Scu(RP��"˦�nkҘzb;6�*��W�/z��cRVNyr�"��2r��Ѣ�6������۽k+;���=�>��xH.�w�������;F���C	:}.��G����T�|O{)B�m�]ᯃ�������%ц�>���mq#�$�:Iv������j��QA��ˉ�ӭ��ڢ�e�3�4:ӗ{a2��=���-j�� a�{���{���0���"������~�����V|(�do�\r��ZÄH(�Ҏ��:H6_Iپs!
@��f�F���=�����s��-�N�0�c͎��qw�Τ�I�	sw!u��f8�m�X��\`��4��Ӈ��GUߋ����O���)�I_B\K<k���v��<e���󢹼��c/WI4��%$��N��A����i���E�('v��zd��c���3�/��=$<��:~gh�l���G�����6=։�2=�
<�I�JІ��߼.������;m�я�=u}G��*'��g�Rx����w߳�|�C�Mr��~+�-g�-A��D�{�W�x0�\Ё�RX������(<C���-{yo�r��K��A�t�TWl,
�n@�t�q�ɭ۾n#���>P5;s�-�nWb�$q�+I�T�@&|���A���
E`��-��"�[�����]d�t[^!�ץ����T~~p���`��᷐c:��D�	�x@��=�����0�[X�B�.uF��2�$Z�g��%͐]dn:Lƹw�?#�t�����%Ub�Q������-�h0��ԍ�p��a���p|h��I:��+k허o�M�|"�:Y�?�Ԉ\hu�o�O��lW�@�љ3�
z
�n�%�=�:����l�$#�*˴�^�q��c��X�Ϻ�,�J�fi�B�!>���|�۷��)ٺ�m��������^�Ї��)ď�~��جz��1p_N��w�4Le�jaԩ�J��C]b�	�(���4��ϐ�U 5<#&��jØ������{j�[(��JOϢ��4#
�u�Q^ �,�s}A�s�HיAD�̞Ndr�Q嬿�0h�)K7�����K/�3YH Y�|)��g��C���P��X�*����a��k�l�]*F�<d��w��/��*< �'k0�-�S(��'�2�Xpg�o�����Q��Z��Z�.��Mb-��������� a��l�-�YTQ�D
��mc����o�k���^�\��޳g�^48-]��{��΀�>�2�N�π�McR�B6nCɛ*�t5*x������İezF��陒>����M�߀X�]&͐LH�o@�`��m�8���C_�8@j��C��RoH�t�6/у�_�o\m�b�[ч��к�o.��e�/�"�r*bI��_�뎁���s�����;�i��
�]`�#A���J/v�F�^*[T5�^�B��E�v��~��+~�˱�Kg��n�����2��/� ܎�+�0T���cn�QV�ZO�:���Z���g+�1D�46�.:]b7�]zrN �_1��h����^f�c�l�x1�*ԿÍmǠ��(y�uЏ��h��a�	�7rO�����*4�{���1e�h�����|�m��zZi��R$����,lV�b-�1�a�zFW�Iy�B q�w��W�el�G'Vط�P��@5�D��+&�.p���V�4G+cŎ���� �V|L�@�l��8�bFV�B��
���� TA��ø�I��i����`�����*�H���${=wq.�h/Q�5�`U���XKB豨�g3�ï�:f�8_/5 	@��B0����8`Gg|&P�c�*��N�dPē��$!bi���#�{	�G>�
xB���Pa��UHCE�t�iF��̪Y�w;M	}˹?��<׌E(�J�a��)o{���4�dz��l]�k�HS;lW��j���sC:�{Þȓ�jPB���ů�y$��lo@�Nj�΁G�iN�9�/��}�Q�tLp�NC"S��&R�ـ�ϰ���ⵆ���\�g�׳��$�G_�ݩ۸:0�o�@Ϣ㠧rRouUK��������*m��D�`��j��C��N�u-�ѧpְz�%6h��D�����<�XA�t3��� wՄZ/�����/���P7���!�n���(�Rp��Cd�w�m�/��E���]E��l������"6VR�2n�a����sǁ�o�p�yǨI���� Mb��h�q[�? e޲�,�M�ԥ�w�������i��?�Y�ݺ+��>[�u��~½��}�U��ZW ���4<�Lw\]��(0d�+���9�Ut����]���h�-m�G�t�Y�C3zl&JV�3����{�弓�Z�!�6��L�}��AS����m~{̵�-C��o�B_�k����d�oޭޮt��/Qkx%�XX�CN��ynD���La�Ҧö�M���w��B�����wV�of�Bx����x5��)����*}��Ɨ���!x���Z%M��-�ǶN󥟪�?�[�[��UҞ��2D����#6!�K����,r�;:į��$+�#�{O]!��(B{�On� �aR �O7/����/"��ٳ??��t+��!ۂ����-5����Ď+	�W_K[��\	d_N�5I����D�D���VWTm���6�3+G3X��>=�D@ ˬ�g)@�Lb/.u'��Rnk�ߴ���U�ǛY��Lx���h+�iq�!����H�?���Y=܅��m�i����YM|?��Ryt�x ���V�5~R�k}�E��q�T����Ib�0��ñ�<���:�
0�w+\����Fgd#@F6�V��P�kHp�3�~��������('DJ�M�5����4 e2:61Q|.�wc�_[h4h�Tj�Q�:��C-�o6`r10c��G��fYFE3=�2&g�.~<�:�A��T���L��	�r�$�����jlX%�k�?fR���W;oX?���(V�\L�$GW���9J�%���5~@y��ZǎfY_�)�L-!��(m��/i��@��m7��p8;�R���@{;����sb-�@@%�ТQ����<,�!r*z��'��되�$�̵>���R�"tj���o.���D�&I��bm��.+~�����.��j����D�/��<�.bd�m���i��Ema�`��F]P�j�rY�BHc�����G������֮^����ζ�\��:�mJw�U�}�˷��C�\������bs��t�/���Y��7I |j�$g���ӿ%�����e�I���8�+Ỵ����]Mb�i�!���u���?TwZ�M�ǟU�U�ihh����ż�;����D�Z[�'���W��̸�}.�e\x�U�܈�:�J���|s,�M0L958S�RB��N|��%�B�S�9B#��@�����å�h��P_���O��Btؾ� d�¸ዏw�
�Y�KsY��';Z����덙v�f��.�88���1�Í���q���L��P]�g S����#�x�ӢS���o\� �Ľ��v�������
�2>\�')�[.$�*�wʞ]�(�?��ڕ�x�5�a^��g1�	?f���w�--)����`z�=�9�qn�0~��F��\ ����0T�-���t��a[Df�J�L���e ��d�!��Y�( "-�����_;��t����t��]�,�� }�=J�E��r�^֒j0\�Gy���yh��7��c:VJ�5^�{�1�{"�p����-D#w3嗁b�j������p�3�x��S n�$���}�S**�I�L�O.�h��Ɗ.�z~�$�p�S;�?.�����B0JM��/�kb��@LX�NRA�w�s+A58�"��ۜ��9��.awS����^�L�<��%S|�{��f�ahBQҮ�Ɲ�����)*���l��C*���lr`�T0^&���ta	D�X0Q��ZG_�j�����= �B���h�v!c���*�P�68�1l�<�(7,��%��\21�x�S6�"�nVh�����K�y�͠���B�T~��eӕ�w��h �"�z�z�˅>��iga�"�%K#�� �R����P���t�v��X�qU�;��,�{ڝ:_2�FL����^<`�igX��&2�Lߧ�u�,�I�|x�0_���I!0Rb�c��)�A��Z�FЅ�/�g������n���OԐ���%�K|zN�:���mޛ5�*C�*��NI)��c�'�\�M ����Λ`ȓlQ����Uᑘ��6�G�y����{]*SJz"ׂ	�^ʡ���\��vR�џ��^Ϭ�N��G.��Vש�V����
+�X�~���t��7Sd�d:�W�r�l-�7~E1(-�%䑜�Od`��=���)QŪv�Ϋj��������.J,���Q]�bq��9k�}��&��c���|��
��~�naY�Xn��DB�o(��F.	P}�����{�lfx��l��X!#� �SK��V�'��Kͺ,����\N�F�-�"C��@�T����k���$�����]�Fj�%�%��f@@��5있�����i�O�ׁ�^��\
�/�E2tmSU����u糧�7P�zd���7�":��=�����\XҜ�ۻ�Ǵ$��gp�Oi�J��/d�����P�63��#��/�%�}[��[�x@�_��� �}�,�m��5 t�B5�Y@��5�(o6F��9��_�Je�v=?��;Rܒyhi�}�*=�)�);�x�h�1v�ZD]?�@ͪ.�}H�È�]W65��~O�+؍��I,�Ӥk|��~a��0|�T�Fp�,����jt0��VM!��vޘG�CJ> �I�a�����k����E�ɩ�\G�вyrl�����]����X'�kkqkz�h��;{	���m���B��IN���L4x����7�&i��d�0�YhTZŔ����+��<�ڀd�D�*@j�P�w��@(�q@����*�	� /;tTOb�(�i|��<
�8z �b�.}_/c�\b�6q�߫~*M��������1��jos&��ZZ��CB��0~��r���eة�ވ��ۡ|Ltc�E8�Ci�q�x|u���PI�zm��\�;����1@fw�@�R�0ɽ��.H���?�42gwі2�R�d��~���=x�1���1�A@��8l�.kS����x��cc�<m
�vd�{���o7ñ�ݞ`%k�Z��7\���j���cWͮE>8Q��	���1z��"!Z/~5�L]�}�N8��T���ꗌ����h?�T��oq{��b��7��������r,3L�k';�"]ʄ����,����w�C��B���բ���=#8�5���.�{�㸀�3�;
��>��lx���J�ze�' 5�h_����0-+e�T�M}����W���Q���|h�I�#
c�ë廙|pq���ՊT�m��u'�ϵ�26�4P�o��@JJH;v^�A�՛�q	4?���!ʈ5Lr݃Y	�����4���o��v���u���8W�j��F��ns��Zb�!MSyň7��5�O<��/�ۅ�,���W���a������RQ��8���Z����=x}_8��Z�kbI>��p�������,�-����dy�ݸ,9���i�D9$T��X� �ϣm��D=�X�
Q1�
�Aa�%h7��J�r�O~
�\�\M�S��J/n����פ�Α�48�������L�����6_�X�nG�&bc���d9(��y�H��le}�Xï�:���!��{�
	A��b�K�p�*��6*p.	�"m�-�%�<ٲܹ&�i�T�<U�c�Vёբ#;�Q�yT���;��!tp�R��h֮N@����9�!���C_ol��r�9�6e7���� ���`�5��1��6:��F�hTU�p#pp��tZ�
'��c28q�|�,Z��z�G�[P�Q�M�E�n�̓	��,u|�����Һ�5���F���	�~�hs��rxѫ�� g������}F�)��L�
�S��Ь���t+�Wџ�=��W�G�����,�ܧ��OE��|"�D����E��c���l��З$6ڤ��fD'H<0����3�~B�[X}�g ���Ǣ����qq�2�u[N.C9<>���7�A��'sK���ʱ�9��"A�L�FzYjv,"#d�wGEsG5����+��������{�5�ݣ٪�]�R �K���6ڣ��7wDk��~�d}�A�W�o#5'{F`���V�Qߕ�c��2@�5���F�0yDY��N5��J5OL�ФQ?�v���p��M�s� �Ț%@�g{3������2��X�&Yɖ��У��6����O��Gd΁jH)�?<Ԗ���胠c�i��h���1G�}�����;�N��㬀�ב7|8�x����C��̂���5)>�W���J!��>�O�QB"��Q�?EF]h��:G����7x�\��Rd�1�RU�zY=��9Q������6˻���g���צ�X�c?䢆�$JȘ��� �� ���?��53���2��n�GQ��~T:~2H(�._Z�U"�U��<�ld��-x����썁�^#��:_d^Q��_8�=������5�r5LJ���Ҹq� �|��6����Ў�l��!�Fi���i����2x��E�#�`��xB�r�:��͝]����R!%��v�M�z�D9K��V��q
�畖a��H'7����$E'�8���2�	p"ڲd97�~�D����	�P�3��_R�^�I)SKn߀w1�(�*>LN�VO)�8�q)POM�ΑܒQoL!�8C�]���T�Q������G7���\�rT�=���]f���/�0�n�A<m2	83�Ar��K9논�����ܨ�[�4&ƾn�����pϲՐ�;S$��TJ}F�-P&�c�/�9�2�w}o�ޒ�o}.���e1>�v[Iz	kJj=���,NY������f[��?��.�cZ��x�6`7|��n�,[cwJ��8��ʇVYgQ��SE�ʠ�v�+��W$c<�''�EI(U�������]c���ge��1�����vi�mJzS�UK�}et�֯�����sٗ�)��������w������z�[V�[V�'6v��P˹xֱ+o���h�~���=n���S{V��eW�����b`���M�3��($�B��ng�M�,cҾ�ׅf�'{&�>-E���Z]�*�C1F�v���@ލ���%�?zT�Lhۻ��=��&��s��L�lC-M@Hw0��nx?D��j���uf�DG=�O�Y�X u�8^���n\���#',��I>kb����m2����ˡ��}*~K)�O�lC.�u��`��G	��ݑ
��č\�@�@�^�YoZ�<O�������ڼ@�"�k��٪���T�m��6�R�����jNk�}�Ua�+*X����.�>��b3�2�vOv��5Ca&�����&xJ��-6��W�����g��⎁k��������ʦ>[f2�����$tȠ��IV�-�Κ�ǚx�tx&O�R�t�ʘ�D���:C���(-1��mŢ�{��sg��@�@�����������6:2�w�ߝ8����h��>�B/X���k���/j�/)�8��c�l&�n��$�9���qJ���&a�)�}�u���5���8�p� p��1�n8O����0d����s$w'�Cdt�a#���S
�fr�#���P�k����Y��k%\&Ʈ��OL���������8��C������]���-J��e��xp�A3�eM��#��;AZ�p���j�㓭���+"ǉt���\�űj��!���|S�́��x�-Y��V��ꚬ���o��A���X7"=j����~O
hE��o���X&Ÿ�a�|IM*6ȫJ��ە�eg�`9+��t̿,q�w�-���!M}���gpb %�d��ԃ�Ƚ�"���2��/5��L�P���#�U�����񕘙4l݄&>�h9`AýCd���,�6:z�S0p7���΁�i���gb���� .��Ig�.Mk��c-F��ɒ�3m}a�����l�f(���L���}~�w�KI�z[ k"�qpe�E�E�'�HQ�H��z�xm=�YSb�|�!7z<Y�Ox)Ե�V�:��l����&���&�LQ�����4č�)���`�Hv���S=$�I! ؚ��n�߄т�<��?���'����\�q଼<�1�$T�!�H���i&�|�.G/�v>봼|qǔ�e��IW�V�r�K(���fi Ȫ-�'��EjLm�y�~=�4���WW�����'c���R�ǟ�-�t'5�}M�B�|3����J0�͌��.W��y��K����C��@6����H�#���i;��u]#fyF��kQ$P�{�j��Vw���
���_�ȉ&PᱛIsz�>�+ �����D	�ͺ�p-W��F%���o��ry�z��A�Y�}��Ac3.��@"�[��f�s��� vU���]]W�D���x�>xn�l�Mp�r��"��BMoz�[�qJH�@$��z�s���I�m����v��=�FŕQV��\�`����YB�3J�^P(�M��Ȼ	���]�Zh_ˌ[~�}��bJ%�����Xo�� �m��[AWDp��$�FVW���o��u����q���,}Gƌ�#�����kj�n&;r��"��(����=P4�@�0�����i���3�fXK�Y���r�O�1���\i��p��\��Z�J�v��3R���L����D��������C��tz��+��o��p�H��,�Y�7_�X�j:�3�sx�����T�y4p�t߬#�Q�w�mT���6H}O)=�Ĵ�Ո�$��������V�,�� UD��i��vH�>ߺÚ+�lA�>�W��ޟf��x����k�=쫡4|0����qU�_,�z(S��:��rm�F�vf��Ii�9�-)`z3�o�[h��OڟD�!6�Ə�Kw/��< g���e`m���!���jn+�hN�J:C㋙�KJD/�E�K?�SN�^ar����piD��*��o�
�5������"��xS�&�0���nzS*�-�^��|��L�$K� �	=~V੸����I)m��)WnS���4yK��w^�)�L?�>*�JT@�P̛x�1E����S�	��\[j�l�Wx_!��5�C���Nza��eS�!�	#�C�2���o��F�Ž�	ޭgze�S��c�2�N���3�!�-�=v��楪�X�������5:��t�!����xq\��*��$��"�5��d:���� E��"9(_Z�����f��&���!���r��K��p^S~�t�!���$��d,�cu	~�I��HWw+�١�����|`�x&��#P�E%��8%�v�{��U#��y�)���Vy���|����l'�ǾE�:��U�<��_Z�;T{k˛�,��,<&F�M���(Z������9�gD
7�ն��Qݕ�4��L�Kk�)A��@�u�v�3ٿ��_ەȬ�!j�`�I�ڧ.��aO�ޜ��2B�e'�׊����c��-d��` ��t��t-pEgOY��yjV�w�V.px��7����\7�	�o:OV6�;�1�R�Cw"�?a��{i�|��6��1Jo/\b�/cӫy�h�j~Q�����Y��:[M���b[e4߂��"zW�qG%�-4HwCPt���@!̡S2�8�&?��_���*9����?�}�̅-h-LL棊}1�d2����j(�2���dH���ȥsB�j�U-��o�ѓd��b����-O�?_Z��ݘ�	 �\mQ��^�������+����q�`�b���<�{ݺ~Ok�ۋ ��l�J��>�G�G�쵍��:��]Y�N�I�<�K"��_�T�J�
	�F)����r��bQ��Cs�#����Ď�Fє���f��@�ql;8[ا��ږ��a���b��$��0R�6�5�Zew�OGTj�9y�p��埶7�Ȁ��`Pa�Cd��B::q�Z��9�wIu[��.w��L9�q�
J�玟�
~��&�{�wǖs^����&�%)�h��#�\������u����V��|����:�lF�.܊�_�`�ʮ�}o��D8�y��EQr-ݒ/��a����V�ה��� ��XTw�C���cC��ΎF�\K�B2O�m4�Q�Z:`KF��v齪��A�$��X}.9ۑ�r.�#a�Q�o���6��0~����5�ހ��^�%����e����v�D�Ԍ(���1����k�^����nз�?�7`{��I{~��@�|�Ub����o�{���f�����	n�u�sX�Mˤ�k������J��W&�{xT���K�9�Hn=Uh}5�Bo
aJR��=����	a�<�Xꏠ�'U7'�p��WY���V��_���lk�Ÿ�t�oz�����4L���V`�*.H���Y��L�,�S�$9�'5����[e��_��Go2��t�	�b�IfUj�h�eA�O8�9�;O�%���K��o	4[����K�0����Ѩ�
��&�[)BF�5x[�*~=h;~��<��er$X�^R�C�GQ��g�*������E���(�IHC�xB����C�J�.і���j5��O��5�Q������{	�'������>X�>%,Y�ncPo���[��c�|��t&<w�K㲄�d��8BA%p�p�?�U�al��8���PޖT_���)��*8�t�F�Q�dI�}]�d��u��L!�R���S�]���bKY��g	X�A�!�-�:�
[	�T�i�;��/>q��n<G����C,\��X޸��� ��8����Ƅn��+9Yq�'���SΟp&@Iڗ'�)	o�1 �=����녟6�f����yC�����G���	~�-ƛ���Yˍ���2�%�Bi�u�Ҡ��Ea�G3��Pd/�f`P�J+�(3�R��0եfX�gM44l����H����c��(���Dٻ�3�+,w6`i����9m��C�0yMg'�����#3��x"2b��\1�m�|F�*��^���'?�����q�W&���g�����D+�RE*���ǔ����.�<���F��n>L�'^��b����5��>���L��{?+ }z�m-�2z��ԐE��s�lz#&����M��<м[��wJ�4�+΋ıU9�1�b6�����%HET���_�I��Ĕc�#���Z�
�������m��i�(-Upƅ��Y���|E��:���0_-�����u��RL/�n�_>�"�S	����y.US��7��;uZ�Ҟ6���r��'wT���3pk,�:�Q[ȗtę�m篷xްS�OL���?��  �r�����+�Zn��$���ݣh��[(��	t�9��t����$/���V�K���n$kښ"P�Ĺɛ�� ���?ls �4�(@�pԃha(raK�խ�>f�Ę� ���Q3R��P|;.^����ߖ�n�,xa�޺�� �1/�7X4�Mpӡ�	�&�r\f @N3�f���&c7���Z��9~,�z�_x8����k�T���#��K��<�5eD�(	�0O��R"E�wo�U��tP�U��R�:|��T8����=X����#��n�X<\�s��YS���pk�Fğx�˛�Q�]j��<����V��ɤ�U��H��=[�|_IC0{v�Ȁ�o�E�9���"�=�e�&�Tt^0�G�h���>�z)�5����n?z�W�V��
��.>ٺ�����մς-�	�%/_�����2��2Ex��IjC�������ݑ�D^�+Z�gQ�M\��o������NP���ƫroD`��D.��|�jv��7�:�i�Fk�gb�k���g�9�?-����z���9������^�hER��'�
��#����R8�(�y��G�Q?��Qk&MQ��l���Z��r�E+�����7����S�h�i+Y���JMH�]ڍ�I����_�2<$�H���3�`�|�N`$f����6���B-�q�+��:���3�Q~�����,������H��;�o9ɒ(��8��yst��i5>	�Ҳ����sT [��&�s�{V8h��(��!ZUߣ;��b>�1)�G�BC��x��5����m�^ѱ�^��OL}f!�$/U}B��I�a�.2M4��لfe-�H�[�(p���S5����5�|�9͉������)��,#8�7���G�mߒ;q����b&4L��hEL���?��9K��3�3��������Z��Eඪ���6�� -��P�T9T����7��\�~�e6���M��7:���s�0�q�\�+���H��Z��<��\8����u+��AT1~\o�i����"r��4i�D<�|V�r��Jݢp��²>=�m�8��m}k��m��=���W�-�rIX��R�H��Y�����Y�D۪j, ����:M�%"�s@5�We�W�
�4�jXh�?T�)� N�h��\����6�S���]�x��)��̟���)"��&bF��D�-9�s�gE��Wi���'+
9P��&i��e ��-o�^�xk�=��-�~Ew�M������ϳֱf�~E��SH?�� �C��1�s���+j��gg�X�TA;�Q:.��4]�� ��H@�Z�xc'�=�*\��oE]�<fY7��y2m_f	%_���I�mlq���Bv���p��qZ�MM'�V���&R��%w.z	NY��z�a��W5?�
:�^n�����ҙp�r�
�nёŋݮ�?���H��5e�zfH#iV�.��%D|�A��X����O�6�g�|�d93^��[A�{31�mhҩ�S�j�u��b*��R�;��Wj�ϰ�ye_ݺd��ͳ���H-���� �J�}
w�� 	I� J����Bٌ���ҹAH�ֿ"�T��p����6��RK8O-�&S·�����@&��[8��~���P��L)*lxPR��		�5(�ߣ1�����	ozB\�MU������~�w�!�Ӛ�4��v��<'���G#@���h�16�"�%ʑ8�<�1��K*�a<���?d~6
���;�2�9��'�ɦh�Ot�*��	�S���<h���=��>3���¢�:f�gGw�W��r�~yML��^�M'����k�A�7�]miva�e�,R7 b�Ax���9.�f�[��͸��ut�䜑	��r�{�m^G���h18�Y����>8i�Kj�m���Fj�y���n����XdO���c���4y�I��o
kL�z����<z��y�G�ڜ�f��ASR�cԏfم�@�K�Z�"F���/ym����T��\`9I���t���(�|	���`OR�����(�e'�kmS8 ]���qd&�#D��^ }��A�(P������%�r�ԭ\�
�P]t��	�2� N���qpa��#���8G�ˊ�����s����}�ց��s	�����^�q@��.̓���K��޿M����r	;�j�� ��!Ô7�&��濢?k���tvZ�`��)c1EU�#?���j:��+�)
+�SM�����wa��XS�ۉ�g��e���J��m�|P�n'��;��]�����h�l���]�hhv,��	�w��Y�o{�L���g%��5�c�����z�=$R8�z	. 6���+�`@����@�GV�PY)���V�ܵ�`x�fUz:�(���i���e�d#AYs\�sÿ�+ڕ0����O�ks�6��KP"��т���+�p8�5"�Ց-��9��+ S��5��[�����抹��k� �J.2�ċ�j���:j�+(�.���&�ܨN���Ÿ��*��^�|�V��I%�?��Cʕ���g �K��Q*��9:1-�a��z�oΙ�7H�������QT�)�X���l�s�������AoM��}�������]�2Ϡ�;�s	@Z���9�_�������r��Y~Q������O˳��GͦokO�v��`�Mg���1��|�9�?�������M:��:z��1����W��|����w~q��ԁ]���Sfі��$�:�Q�<L2[�� �)���npn�Kx{Е~���ۂز\�`�k�ElE��N���g
'�
y�����Z�W
�Ӑ��a`_�p>n^Dx�����Ct�s�3S�1y��h��Db)���K�2���CX�<��ߓ�Q�׳2�4�����	P��'=��i�1m	n�5v�8�������D���������54NO�������4|y�,\��k��.�hT��Рi4:`� v�kق�y�f�c؏���#�I>�7�l������*�h�R�[?y¡W0k��CA�H��M�D�[1��~A�aO��NԞ2��U��K�i �1���h���p�8��[�^�3ͩ��iP������c���74�FWnUcp�hA���ÿwG=�Z�#.�2�*z%}�|~3�qz +Xޤ�����f١���4~���XSG:�.@t1HV�nK�����Pέe&<&y�(0����h��Wߜ�k��X�bM�p#�=|��19�c����1 �R��J�zs���N��9����l�������?���F>Z�Sc�Xܼ��9�սd�P�B��j$((� PTYh��{HpA�ݜ^.���xn"��lb*8���O�����Ǌ"�-R,4���D��i�NM����~��5��&�HXY����4τ�Ͼ�f5�fa�V/3T���ZG�\��|th���
!8���8Ўúݑ'���b������ �����`�M�Jt�p0>8+��i�0�i�Q�E�F�hï�ɨ��1mw�\n#}d�[�ڪ�� J�u�c4$�ٱ=�S~d=�u���Z�FrJ|"��j΂�)Y���ə�K"b��A�����mcl��������S��	!�0�_]��
�k�E�dI��i����!d`�E�;�.%���#��sz�TW��{����E���b
4/e��q��l���s�?.[�����f��-וw��f�ɰ��oK�J�3�c���1���W���@ʨN��BY��.���ugc�p���a���U�KR�M�,t������Ѯ.�ʅ(���Ȩ�c㼃&�M�������m��9.=q�] HJGQc-����f�6T[�$�jo�(�'��p/�pȬCO�s�^}锫{�-�;��ӯ��f�\q׏�s�o��H#�,���
6:^Ajҧ<���5tA��Z�>�	Aa娸N䇔@9�����mN�=�W?8!}�7n��#_h�W����WFj�0wS�9�%Gh��Jd`�[�}kF��Y�����|���=X�w�&����3�+��jn]l!_P�w�f���d(|Q!^o/�1�*Ƅ�xi�K�SZ�vo.��x�k��u��=�i���/iK�`K��~�Vd�9�6T"O�&��5N9Y6R ��p8��xsӉ����"��UV檤s��ؐdS���q/�p�JL���8m���\GAj��d]O��U.���{�Ji�I �� �3�$O�o��qg(2I���3/���d�eG��8x�Z�.B8A��(����~�Ǚ���������O?�@�k���$f�����IM�|F��HGr�W��S�m�C�4HD?��:� ������)�֏Ñ��,�� ����X� )�g8����s!ڏ��N�s�K�/\@�|7\�N:]H�
t�p�ZfY�~��M�
��r��i��⍤�%�p�`CU��߮���jW;�Y!ԏXd�4�;9�#���D�r���ώ�y�-��ViZ�G�����7��U\��t�hx
���4"����&�����2z�Kj07I����O1��Ȃ�M�D�f+ư��_""�n^�u�)g�u���K�i[BM��͔d��F��[}��V&� �f.��-3[�֖���?>R��|2��kR�2�ie�U��8D�ͣ� ��o| KQK�	يԏq{�Ó��~$6��n�9{;�tB�7�N�D)Wb���w������� 
s���D�u2]}M���- 9⎵�Y������.��K�kB�>2��*l��_OzJ_a��$[�.(:�g��$�c���Cc�(7Wӯ�Y�`���Ee��E�Q6���wLF�Z����ȉ���Ō����}��|�{Zw����]������\¥_�j���&�e���v���n0Ll3�r=� ��ú��+�W
����f���h�����瑄�G�Ou�&T�8;�+#N7u��T`����d�V�;��p��D�^�4e��Ґ����N���إ~�YŸ�T,RD��	�T�5�Y�ÅU�ʝ�mM ��-�K>��	���Վ�)̆���W�s?�%k ��&I���	���#��䓋���v�P�H�SauBQq-���L�A�]�@x͟�]7BRI��pkq����;�h ڼ3SHj����0�4��� �a^3��Yi$��'� z�6�S�r��X'�������������4��NX��US��qÿ�k7�T`�P�� ��"�ʋ����4�`6�2�uf:%��C�zK
�f����������L<�Y�X�1ߟ�74����4�elκv��@ށr�>��pv��B�f�!@��
�}]��?���Y�&�]��u:��C;Y}||�ph�<i*�<�������u�q�"�`���Q
��`>42����v{����\_f���bR&�����tHj����@Gc8������m-m������e�GI��Y�Ѓ�ݣeϼ����c�4�b���u��y}s�4n'������V춋�L�e��"��Xx��)&)��\x�ˉ>�B$e�N�$�[��)mt�t~�2y"\aTB�1�{�M��C��j80��)��+�t"��(n�)�Rt��g>Xo%L�k�)g���VY�Um����l
�.��T7~�x���B��i�~��4	$i���)��>	A���2��<GS�8�c�'ϟ�L�sʱ��ೇ�"l��q�Ŧ>��?��R	�g��M�"s�����@E�R��Gv3��1�~��/P"ߺ�_��1����˥�#�_�-����}3��-����&�ҫ��sX��߯��2�19�v���Hj�X���yڊ��(��7V̍3�}ì`�2c�ϻ���,\Ā�� ΟT5�)p�۔<;V�f�A�������ܗv�i�'�U|}�*��M��;�M�kp���GS&򲓈"A�PpTI���L9��.)57x��l�=WW�Na�M�]'��<3�@[�����KS���y����"�^�[��=�%	����#�u���8n�G6�K�*m���w��� oZ��7_ws���׺�\Ҩv�������&���z� ��@x��ER�3j4W6j��81! m�*�6�&�_���ᙻX@:_�x�S�����.r�A���p�[�4�؞� ��h�tў]]�q������։���j�[)����{� ��V;��s5�(%s�MA)��8���B��%KN���MҝN�a�BՇ��&Jσ0mv:�}'6-!���w������q����&L�tlg�I7.w{z��oM!҂Y��.� `�O?1�D�1)Bf���Ң����^�JX>�,��{����t���W;���N���D8��!3S�
 }��JGܾ�\���nK,^_�r �\�J���N�N�8���s*��+e��X�j���'>ua�Z���3�_(��T`���45/�wH���M�%��yl�������xA��1s��u���>�o-�
X��Hw�����ז������.$��aƵ���Q4L��zyv��q$Ә@���lD�8cYiR�ILv�Y��������*�e���+��m�ϡbw#r�D�� �2R  �����Ds�֛����_ᐏ�H����V:���++ r�V��ZZ�=x��<l���4����7�;�I�����d���E����jV�6+��8�I��^�(�r���ŇK�7����Jd�@���8f�k)�Ҷ)��������4Kq�g�'?r���}���N�M����D�S�~t�?Q��f��`�T�����-���ݺ(��Z0e���B5��LoVsr+P�Fk�7T������*@�?V�5�u_�?��.L"W�U*���;�����o��@����t�ވR��.�5PRh!'�'#�9�߬�`�G߫�~�����ɂ�j�8t�%�j>4�b�;��*�fMY����a$�\�[W���(y�;kۘ�<"ы<�m	dsl�|�#,��6�N��]i�Ɯ$(�Β����b5AB�������7W	�j��S<�8ux��z��&�7~���O^��ç�ng�V$�(}����߹�С�z0[Y���ў؋�ˏ%e����/\�hyzڿΔ�M�sns�ޢ�ۢ��E�Ȁ�y��<4��zT�^c�^$|��3\��$���t�hdJj�q�hf'=Z�l��������*x?ҎZl�yy-�m�ߘD�c��6)���,R�	��㇝��V3ULc;{7�5��Q�.�x�+��tr����r�\� H�C���+�����
e�G�Jl'�#��c��;U��I����im�
�?�a:�̉����-QI��T�K�{��ǲ	]�t�i؇7���j٦��*e"�����Ѧ���������g�u�D�����W7Qs�;�`{,_�*�6�c����L����U�&�9�2�5�䔰��$��X��{��r���t�M�0��U��q� 0�r����ǋ���N���Bn��G%���y�P/��?���i$i2�?�+H�V6A���z��i�D�S`���ľ�c5-Mw��a��O��i4�s�4�+gk�.�_m#3W�5&���H�n�]�G����Id���&k3x^�H_@Ͼ�<Ɨ)�=mC�}���%���H�$B�'=Tw"�	�\�����癋j�5��2#�th��o�2Ή�UZ��)2#�S\�|Ua����qJ�5eu4�M��b�/����������R�lu5��mz[�ͣ�ux��������o��Z2���n�P�\�p6+⡖��y����B�>���!�L}�FP�0�F��Bz�6~�<>zGB��(�:r���Q7��3������^�,z�
=^�{zˀ�!�NIJ|���U�W��F�M�l2�:q�W�%6���e�pg���}���ȼ��e�+&���fȹO?�sk�4;5|�(�n�G��x��8i}	6�c��Ju�3�4���:�?5�4~��\m�?26��o�n>���2i��׋fs�꺖��C#d5��cZ���R���1���'��Н0?n�V܊�nN)zN�`U0�..av����%��)���8��F�Y�5B&=F�U@���K_��0�/s|t���Z��*Rg$�˺��<9�
4�n/N�M;g�C��f�|`�R_i�/���c��-S�&�LxҒ�p�������ۙoF>o~���t��Z	����Uw��lQ�N�䟐5�P���4t�b���� �`= ���iU[Dj%�g϶\F#�˪�q?y�(��_�<�(��3�E*۾��Mqq@U��jP�k����X&L��EPA�x9]��~�(�����Ϫ��z2�ʤ���m���pצ;\BE!6
����ݨ���K�B����@��j�>{Uh�G�2����t�9�e�(-\�������d��*�ɥşaD�
�G<X������uj�f�I_��.�?�	�z&M�qj}���Fgxw�� ŗU+�_u��xG��_�eJ��XJ�����d�[`h:#�.0�����A�V��ʅ��Tm;��J�i����"H܃��+�}>p�:�A�Ӊ�!8��̞�@�S��G߽M��`4N+�9T�����>�\��qq���J��71ʹ�].��gGI�z����᜽���f��m��g؁&u����/���Uk��𺉄\�)?�5&b\�oO6�-�C�D����5e��_���f�!�Y9�����W������1�ݖ��x�W7̼�ӄ_Xg�u��{������ъ�$2g�I8f���nX��z��I������4�n����F�C� 街���g?pv6�1F�TR�H�04�����JT��� ��7#�P)���ӈ����&�[3O>�����(bU���aE�)����+�z�llW��4�\�T#bE�M�t��0�PBO�	f*��/H��L�!j2�6[il������7�f)
oJ�Uꈾ�d�4!�-':��n���p��h��_�^,�Q��l0��
(��ux���Y���"븍��f��[�{̔Y�م	�%�7R�IQ�-�"S,�{ǜܡ��a�뤆A���r�� �K��&�;��ʄPUrw��DX�9�M�b�XZ;:�I�\���\݅�S�<�z�^�S�8��U����kX1������A�a��?�.+[�|����d\����B(!�exv �ʘn!��Gu�{���	�Ӈ3d;�-�4����>R��Y"�����C�yM9�������}U�b� R�^���o�\�L�#8FP�ԟ�Qt���a��Rt�4d������7b�%��׺1˔2̲�N7�d���O��"Z[��7�5���Nu���Z5� ��.9ޤ2`�K�C�\X��t�_�1!�1BM�y�lL~`2E^	�cڗ��K��Q�vn(e��ߙr�y�J7T��x�U�7$�Q/�����LZ�O��M�摦LU��-갳�Z��}!u��B�ޒ��D��X�m%�2A���BQ�b�̲O�NHث  _�4���x��9C�D�O�(|�<'+C0�iw`����>,�]џ
l�䰋�6�͙���(ѱ�Fyg��rEk���P7�!�]'��rñhd'�cҏ�s�1�$lx�N�Dĩ;s����ky,������6�ه�L��8y=Ϙ��u�E!H`-$���-CZ�Q��_��`ܦ&Ŧ�(�{_c}�����㋕+(�d�$��HQP�|�䲻/��Yc q>HV��k���d�գ�"i�z�7<�d��S5`rC4!��F����V���A��=؞��kϸqf�z	 ��c��n���*;��z*lZb�׏s�=����Y�RI�sap�߈3�X�T�r>���J��c�-#��6=�r�r֤mmOE�,����i�,��DH�����M��1.���i����"��q~�J%�ɿ����"�d��m,�q�I��߮u.��od��g �Q�?WY����)Nu����5n���
�L����S�1'�g�XX��eĿM�Ԁ�腁����y���U;_U�4�`4�j��G���N�H��M��t4���j��Pt����Sy+m6r�dw�^�J�qR����\�M���ߦlsQ����9�p,QJ�Rum;�f�_�Ξ��l�K_E�GB!���Ί�J�2����	jL� ؠ̨nE�n;�v�3U+�V��h��L���+��ú���3��,�Sՠ�gˌ�p����"�kbv�੷��u���&��T�ώE��3�����Μ��W��x�2����l�8�7t���	�&VP����Y%���%F���eҤ�'��?=�i�
�$V��T���貅���&ƌ<<.�x1�1)�j<+�!��rER���z���[ !zבFp�#[���%�e� >��SVz1���$�DHv[D��G���8����+j�ǆ:|˶[��:u;��#�7�){��**�i��I#C�ٲrI�%��O��i�́0q����2���MO&���\��"j�L\E%O2c>͔�.����f6�Y�G��������֩O:���c-އ�Q�fN��&Ia�,`Z�9ƶY�|���ANC�'�ך-@㯏�'�k��h�蘚Rr��� V��+� �Wς�[lr�֔!؆�]���{���,�&2����O��rJ�-�:�w�kaO&��۹�(���{�cCb�@T����U����*.P�@r�f�+��h�DU�)V�ʆ`���X�(@]JRsjl-J��IM�w�, ��u{MK�}iZ�y�/�p��V��v�$mթ��c�v�`���6��=@ƽ�tW�R���l�a*J��MW)8�Ju�M
�7'�� �z��w��WQF�KH����M��r+�ϔ��	��OF35d�S �;M|�(�^�,j3�4�i������W����6�DG�=t�tS�����̐�[oЈ�A�݈���+]�`_t$M��6���b�"�ܗ���Vyu�"�%��w��_f�N�\q�F����\��8�~ � �G)3������P͛��8��x���n�;P^}H��0&lR��Δ���I�+@1[���_q+��#eD���FUM8�ݝ(�;˽\���\���:��v�H�=�Z�����50�0��n�$R����s\�6�E��Z�ω�|��a�)� j��0�.1.���e��^'vx�	nU=�|�E7e&���sU��.)-<�
N�ƎԤ��P�.�ôew�ܪYv�T���<%Xm���������wW��g[�k�:<�O����}�o���@8EOb'���#�S�Ug�0;�ﾑ�,]~��EI�X�tm�«B�<������:1��V&�iC��_��`7m�����#^������b����,uI'C�&p�e�.���&�q�C�L���fba��aۣ�ϖ^�A� �����ws{$��q+��Bղ�F�5LښC���u]벖����y��t�X��5X 켵�5���Gv_nf��ႌ�W�".uYO0G�l<���W�>KEI�H�e8�����Y��B�G1������4x��i��*hV7�q?[� P	|�CD��W�����T�z��Hgrq˹7�d�
������?uش�����X"�n�rF�
��K���oGf����EGN�9�7Z6d�AB�+H����d	9���sẒ�5�*�P�i�/4O��9S�Po㨹�5��Q-N+;ض?�`�<��ț֒#P��	B�H�:�����Bϫ��]�U�!�H �~䦜����+�� ����kU��︯���y�����8 	Z��J~�r	�U�Q%�	m�r�G�5ܲ�-(嵯GpA^C��(�~�GѲ�QW�K�J�:rR�'���{ǅ�x�s6D�q�����Ϋ�����\�q̵�w�����"D�S�F���R�}Hq��}��y�r�5�c�}��è /fE�#.��y:J��e�]��h��%����\���'c��O��
TL}� W�����O��|:�jUY|�5l�՗Vs��8��}��l�F8��H'e��n����ɍ�w�ߋRh�b1~��I�Xk܋��O�Ԗ�	�=ZJ[2M�34BƖAOF�ΚK���y�:�1�'�^"l�Z���q�\Fyߙ6.���dp�ޖ|�VK���� v�fȦ}��HXƹ�ⴛN}���z�
Ue�z94�|F[���J5�R6�*s�s�#b�\hr5���
���¹7#�L��q/89�����nM]BBh����h}ݶ��e��S���|
�]�Z�U�j�l�YdPr̐��'��@��<`������ߎ��'{����+��U��m�W݃�r�-�D1�	<G
��c�*4iƿ�\|����f�������`Q�w�����5%�<�`�i�N��{�*'`b���oÑ(~3�<�頄��$��R�D�[��ρ/1dT��_�r��q�ɲ�)��^��	O��.��0�(4�u�B�b��8O턗K/�)q\��:_۶��>P$��>{���18Q��nS���W�Y0i���h�~>k㳫�QK�HԒ���X�@3���l�J�+[��agf��Y܅���7��d)��4ҴtpZ4�� �>o��=�f�؋���������]]���ծ+Q��f����Vd!�4K6t,��)��G�T���*��,��s�?�$���{(�:�,�۟�%�'f�&��o�]4�͌�_�&Jؤ�Yc�����D�[�����␶ �E(^�w
`���������*�}����5��4)�� G���o<ue���ECc+��}�.tp"�iR6=x�� ���.����p�#:*�k<'�e��x�&�,� �ltO�Uϔ8��k�H��A�ꤐ�qސ���q)�N����: 1�<�{�Qll?���?@Eh?���-yIh���1�U����i[W��FXS�Y=D�M"��+Ibz�?3-.Oi�>ޣm�D�"���L�Ί�	�����yb.M+Y%�r������j�=|���HG�����7e^iS?f[��q� ���i �i��(�p���Ű�p�:ns~[z����H��c�>D�i�,�d�1�0*Ֆ},���<��~���e- �o �8�n�\�^c��T�=C���3���u�u�;R�X����.-��y�p�����HB}��~��,��!,�V���3l/j���L���lzn��~b��3i嬽k.s���=`)^�=6��B227@��i�]�' �d
�Uò�0Gns����ȴRqMJ19\B�%��$��9���F\��W�+��$����rwy%ၘ��'���ጉ�A���o��Q��b\���/x)rI/��������Υ��'9Ev��H�M���7��g�վ;{���@�2Z$�);(љK�	֯4�~��.t�x�G���*$�wԏ�4�Z�2��b!7kA~)"s�gq9���Dwe���-}�J��f��$�����(j��b��}rz�רj�4t�p('�)}�~UWIt�ms��/��99!)LE�&sA�������;�3ݟ�E���"���=���ͭ+F�E�WVX5�f�"����<�3�/x}_y�g}:�Y���op�Hs�߲�#6*)hv'Œ��}�����ZN4��Z ~���eR]lF��G_�U��x|uL/����Ux@��e����ش��g=�~iȯ�&�Z��Y���~�j<�ZBHF��������ƤFJK� w=iQ��;��#:��=� _J��os�?�� �<�y�#��# Y9��"t k�:o9$vC޴g�lH�j:��$���v�#�2�*����t�Ṥ�i5���g��j%E*%A����x�����+��$K����Z}7mk���U�������QW�[& ��}r2��`��T����;�:__����PE���&�r����y��������V/�	�T>�zb����5���F�~Ƅ�t��N�Hd<�mȡ�My��e:������a��sk��!%Bn��a<����#3;gv���]�m���uد/��,�W"�E��Z7�?�A+��9���|�w ��ֱ�@a�T�h���{c���:C@pbo ��c�
V����kP�m���=����=RU�c N�)����փ�kY��(?&�&�4����y�S���0���?(sV=��Ep���c��/o�����۪��@o8���m������>�W�����$l!�4'ڇ��?���l�w�7�S��Z�|_,����VH���zE�u��&Cg 0a֠R����jS<�fS�����J�����I�C�'�!=�/*���1qY)��G��PF��}�8��U�r�y����g��@�F��o�銎�� Gms}��"|s3=1�c����F{�.�$�>��Ϩ���]�����c��܅ųQ\�>w�@BȌ��Y�F�;��*�9y�����ؑ+|6	�h�ڞX�>wz>���=��e�y�a^�о좁��.ĂҥI����§���*�L������Ǚ�L�rJs��	��ԏ�d&/ "�Ꙩ|+�
��{c�p�{u�,2�E�uy�M5cH�Ѝ�7�z��ғ)?�h� �yM$:��x�{b)P�(�J���Kb=��Wfq��H�_j������%����:���"����%9p'�X���VE_r�}Ŗ�2qE N����/�I#	i'����Q��f��b���d6E�Y��>^�dv�"�ϳ��q�k�/}�һOe�S��yg��cX�YiB��m�y�t�X>2t`�l�����;��!��Q�gP�*���
�P�|��T����Ȁ5��n'��o�;��AP�gB]�VD�n�9NJ5�F.����s�+�f�X��Wܒ/���ˡ>���μ�$
d*�����G�Jˤ�`�U'E�2d�|��w�e�޽��C�e=a\Ci�H��Ug���tƩ����Bs/��Rh�P�rc&��k����u<SZ�%��7��c{�)�ߛ�E3_�6ݜ�O��}xė��re��j#�c�)����E�_q����ao���k��:���i�<|�ա�u��'����w��V�KV��uD}듅����(��x��c<){}ʋ��w�"�~�X�������8��ڤN*�K�'q�b(j-�GV�8��F���M���
��I@���)�x	e3��6T<���~'D��+���*�g2��P2<O&�!��h���ЌF0���5B���R�🻄S+ה�����T�P��f
�]�a��Sb��\wj��ħ�b������A��+ja��Z<�9V�"\���Vu�����}W�&���V-������m�,D-fr�1|$�3��\\��._�qەL��4O�AW�}���|9�>y�wѾf����܎���`:�Ʈ�v�1�I���1<��o�甇���|*?ܲ���j��w�OI��c�\��&�Pߺ(�k�0���'�`aRY�'�r�E��t�+�V��V�<��.�5ň�Ŋp �3���Z�	�ӷ?'��hA�Q��<�ş�:�� ښ���Lgw��j�%�]���&��`�:1�9�����&�P�<�R�z��v���=�JBxT�ۅ�-������S���=�f�L���l�x�e�� N��s�3
p:tp˶�����MF�/D�ݱ/"�S��l��]7M��1�6�����)4�\�
T*�XJG����*�����ir{߳���k���,���"Ry�b_��_ �Ȅ�k���Zo}O�P�R��{ռ��a|�"�{U��]k2��*�}`ԦTV~�D�{n�]Uh(�Z#0I
ixx�:�)����sи}P.e�Uw÷�ݠ%���2=���2. ;۴7[Qן�&���!̊������Z��J=���y����U�,"!�Ȼ�͜f�#L��9C�1�E|���I��H��h:*R���:��=&)�+D������O?�ξ9�^��7O���A�u!%��eyK�i_(li�x�� Uo����h##���Ǻ�����;�(��R甃Ƚm����kF������t��J�Hl\�y��)43�צ�� ��J�N��n��TJ��Ԏ2'\�K��`�������j�)� C��	p����ă�^�ǜ��nݘx�Yj ��_۬[�����e����$H�Cʞ��&���k�q�̓�ʳQq��Y$�#[X�R�α�~�s-�����CVC������>��V|a��kq���͹p�M.v�O�h|ӣ���j�p��׮R� �|�>=u,EN��>��c(n?�#�D�!P H�m�0.-��'�(��1��c� "TOe|��m_����V�5Yԣ��3o��qf+5�1�~��E�7�g��p��B�� �2S�H��o���D��ITD��L�=��_���h�q�]1}�Q`N�=j�ᜩl7zx�)ȷ������k���Pj��`�)���$h���O�9O��Bu�0rh���[LH���R�J��|3p�W�J��c֢���gO�r�i�pQ�.���������=1 rה�����
0+��{>(cI�1�q5�9p�A�U��iRm#�(�NGJ;6%�j,�%��짰�;@S�0���uvyS��SIg'�B`��'
��]�g���f�n��O�9o��I�r꿒�х�L,�4�c�+Sk��$���4#9�sLQ�2͂���Ay(1^j
1=iA���>������I��Rc�a�l����F�(ϟ��8N�LC���~����-̠�g�m�<��M:7&9�l 	�b���s����U�@�7�i?�ϔf��A���P��J��_V5P�MKDAv�Xq{��R��\�kd8F��ݫ��˛��:�)Vvf�6��;�i��GU����;
�j4���6"�p�*�}��^%��C��h���� c�p����2���A;E��}3�Z[�`�̡�$��4LT�������x,6�;
�BL>�u�ӯ>w��A�<�A��=d�a(i����eQU�'����2;�]� �{;^�R�SV���m��#
�`|T&z�R��!�=�d|�-�l����G�����ii,2����,�h���xÅ1Y�I�Zι���vd?��ϵ� ���k��EСo0��C���%Bw�[���a������xK��|�f�����T\׭�%C�R�N�V�8�+d����E(N�����]����Y8��1\��K���!���iZႁ�R�EU:o �r��K[����h����;��@��f2 �6U�|Ϲ�u}"��4%��A;��	�?�蒶��?�5�ԕ��ㄏ�6;
����mi�N�y�r��\�
"��I�&/�J�������T����Q��K%�{��q`=2�)+���T����aNGЈ��կ8L�h:�� {m�/�*]]�A��{V;?ۄl���(��Z��I+�rk��̅�=tȌ���26T��c8 ŵT�:?�KB��7E�����۪�Yy����k�)���J��������z��v���p{�69H��O�H=���!_TL��J����;��eaŠغ�1�n�8�|R<H�p�qD��w�JΡo*L��2\��Z�S�hۧ��@�( ?��罤R� pi޺�7W��b89�uM��#���G��]���eҍ.�x�c��&5�3��i�L��R3~�?��Y8���E���1F��J��'�Ǎ��.��l�դ9����[S̽P�z�����<5o&Ĥ���R0�<�-�q�!:W�^���06�+2�_{:�B�A=�bO|��G\S4���ڣ$���O��-����7	[��赈�_tS�ݠ�!.���z�"���J3���[lB�R�uR��N�ß%%�t.:TӰ��B�Zop����6�x��r.3��d&e��%`������[�=�&���`��r�"�*~"0�a�R,kԇ#Uz05��$�����z�M���tP���Lz�R��#=��dt����*$*F^�NT|/�E�D7�_ł�zI� ��9�a�8<?���q�D.��&^}��h���@^!9��բ�Ux�y��T�"���d�qb�c�=����C�������o�[[e��#c�~�|]vl��豊G�:P+l�A��^�o!>x3���9��^b��_��nm���kH�%r�魐;.�5׉���9�=؞���OXZ-+-M��;�«l����O#��[��3F;�.������U$�p�Ot�<����k-���a��nP�c���
_nf��y�Xfq�=6�<+����ve�>��Ά�_w���T~(�ޒF�gZ�eҵ ���;aۨ�o�vb�^ �[�1�Mʜ76�9	�l��V�^�9L����ۅ�Y̕_:�GCU,X��<&u���N�I�RF��N�������'8�x���� �L�n��n
g�ɱ����oݦ����v)P�ȓ{�qD���5?;r#}��s��/�&�~�c<sw�mUpX�A3�+���)l"�#n�wx�Ȇ|� :�PT ���$7t�xc����]�%�}�Aq���q����F�%�6��ѣq���VW����E�(i2��&�"姛87x�)�d�A{!W���K�u'l��zR��q���yL_�J*("��,��Nk�EB\���a��BX�LC(Ͱk���T����FҁO��w!�ui����-��3��{P�w�sV�XHBamWZ������Zv���FL"Y��M=�.����4)�r>�P�<�c�k,��_FC�(��)N�M���t��G2������n�li#2�س�e	y� ����n�W]~�3����D�
�,А�i����u.��{6S׿��l��Nu[�����F�������W���jo�j��w�URo���oe����3�s�3NN��zk�Ƹ���b x����n���ד~�T��C��p7��p�3�ᰧ�aeÒ�qr�F5�p�z�G�v�=���˫.�iM�G(���1G�z%Qx��<��G����"t���A3�_TՏ&�����)^a�j�=��Vu7�u�_� �y�bmvLQ�ԫ�}w��B0���q�vM큡��	3��C>s5�|��W|���t](�V�6�t4�{��ǡ�	��C�8���#;�؄t�UM���hn��qi�a�Kv��d��£_Dzފ�{��y�3V��W��#�J�_s]P=>�j+�g�:�hY#��-�YP� t����סVjo�2��ܩ�׹��n��7��(��c`{����(��i5H�)���3�t-~+�=Ţ��iq/�Z�5v���4�<�3��.o7��*c���m�1"�B26�Ei����Ӂ��̌qcS� G�
6�"f�T���z�тo�A7�_bR*&^���/�!�)��+�·�S�jg\H �F�O��P�!z���U�]:� \q����o�I0���~�b�Hh�r��R���yٲ��z��9��/�����Q����}����4m�����	+��D��#`{����	���7Ft�{$��+X��UO�/�u%��o"���c�*���ܑV�[�o�Q��P��9N��8`Tʇ�+Sv""��e�V���{!3H_ƃv���#𚑆����B��|e�Рف�^?t�L�'�ۚW��f���g���ƫ�Xρ�$��Ur:��&�l���l$�ь��Xx��ՀYl��r&b�b��Ǚk�M�UHm���\`(ÚE>�>a�Ԇ���1�7�$���r�����7B�(�g1asS����O�"p�����CE���Sr	݈���
�}y��L\��:m"@+B�Ǹ���=�s�EF�^����K��O�~0a>g�(�
R|���a����8�ЗWXVuFUf�դ�wν�M:�;]0߮^�ы/�þ�; 7n��i�_�oow��8ͰX��չK� ���n��3b�m2�uio�$� ���������hC!�sr�x�����/�5⦘ ����o��Dp�����_&P��A8sV�7�G�P��S���l�U�*s
�P�!�a'�T�se�ς'�=D�1�_�V�����&�@?��������G��<'A����^fU[����Uwy��'!�e���g��i.��4*�3���ha�oׄotx<g�_�L]�@�Ֆ�t�)K١�{�X��w�0������1[�X�w���eAz�`�u�B5���h�ު�t��3	CF[���KÒ�9`����e�1!��w֬�sB+�7~��&�=�WZ�k�$�͵�o]��+\^�&�ď��`)���d��MK�ۡD��"fǮ2��#����J�PE����IU�#���Bu�ў����k��K1�4AV\�;�_�/���N��<��3���.��'Ѻ��Q��E�ޚ�y򰕏
A��-�j~#�D�g���<z��q���@u^9		�q�w�����®p� ���w��~JS$��vr����b���נq��% ���=�m�~"�#/�r�5k�opA^��t5��kM�e�h��ܞ~TZ�?Z�(��һ�ˌ1?��M�fgo�m��h]������A�����6 j�������b򁴁h%M�W�i�-3N����ȓ�w��l�bsf_Ԅz^+���0jJ�z���+�K�	[�̓/x����>j�P� ��RfI�1t��偨v��Z�Ӗ�h<���E��������1^`w�3Q���,��kq�^߿��ҩ�r�8�'�A�#@�G�2������ߔ�E��G�|2&:�0��C�8�=t�3Y*_��p�Z�C�]��Wmt�#�À��XĆbNZ�#�b]8�"�Z�-���8-��� ���DတWk4JxR�辶��N��Ή��I.M��ؼ�ݹ�T�t��-�l�e�AK�M��d�+?jRo�~���ʰ�Y��>W�Ǐ��1x�G���7����[��̦Of��"%[2��Z�|��i��LE�KD�)��Ge���#���G�ƶR�c���{IU��0!�H�]�;g������aҐ(�R'�\����60V���W��`�n�>��!�6.ꝡ'��K!dB`�*be�*��.	�v���XS�n��P������� �O
GS#�t�/�>��l�lr��&�{�+tKY� �E����Q����[���j�QŚ+].�d��!᫱(�Ț�٠\��#�S'��Q�'��Ǌ����m�4�H���ސdby������;P�SV�Ѥ5��q�� �`�Z��ss�@�����e���)FW|�NQ&i��,G�T~^�"����ʳV�5��cv☆[&�Cג�CM�a����{�o�=T^�!Y=٪ ���1�t�1Mk�ڨ�]��'���j?��wXd����Dn�,��[V�FWJ#��ΌE��t�^}'<x!o���Qb�o,B�jKkM�ek�n7�Vk?��h��W� ��j��P���������e^�ˀ��:Rue ]x���(��7�y^շi]���ᤊA>I�?�	�<��dH�UH�v-!���`U?(��Ii�8�{<G�8o
O�k��Ӷ��3sZe,��i챨:B�zL�F�~��v�buXP7����t	�r�Y?������q��7�r��/}��]�~��ʉ�ؗu�:n�� �*������[�#Ɓ��Pg|3(�Z1U׹,��;;Z3Q?P� 9��#�Y�-_�{_Nژ�V��/��(��ݤw���^Ī?�ڈ��N���4�'����j�������u����']]?�<���?�L��-�%J=x�
�v�fMׇzd*��p�V@����1���d熇o;�kB�	y��/�w��~�&��~{�]C�oo>y;�/�S� �j��$_���b�K[5���׋,���?##}��/:f\�vQR��z�)Y��*�OA�$�8@���T���SY�rdȅ��������?"���4�#S�o�T>�S�0�G�>�})�rj�1���9��]c��;|T���	@d���D~}
���/c�eL�r6B&��t}����ѧ����#B:om��)C��[8U"J���� :���!1z��iʭ�P�gD�)ο�+��qt��+�tad��3��ܠ�8��*?�E����B�h8���_'���=}�M�ˬ�G��zc��UX� d��KD�qO�������;��$~��)�T���5���@�/�0��r�T����z�=/��N��r3�ˬP�P��n����U`�7�s��m�T�"�^�ې*ԧwn��`�����'�-�C��邌?p��i;�m-%�*֐p����W�);G��G����|FN��6���<n�G:s����A�͆I��|Į�j,�bc9�WIΒy�.)��S��K��]�n%ϛh�@����9�[�/Ц㱌F�)�}Ghb�G�)�>_G�#�/�fxt�̕���!�O�����`��k$����0!�O�"���:+L�ƿ
��{Y��9����ML��� wT���f�˴�f3�w����Dj\��of�M{����Z�6=f�>YB��Q@}u=��Z�l��CQj�f]�	KtCG�i#�v� d�����A|����.��b�HrFa�^Ð^�:�ԙF�,V�]�B�Bx�ϓҙ��6
#E�0#bsU�_\m�Kfe��9��$)��r��H*���l�m��2��w���7r�Y�ѻ���)ޝy�b�e�,��_y-�/�����h�_���,8��<WNV����,�jqo��[�X��e���b�-�I�(zvd�v<�M�B���I1��(���c�����Av�c��*�+(J
[���dw:γ_�Jqfg�
��1��z�F#a?5+�}���;
��OT$2�Iק�Q��kir̢+g'�B��F~g�`��׊P�I홶�+����UjJ���v_\!�4O�DbxByշ'H8�`���2����||r�Q�I5YlV�J�X�N���m�yK�q~��^4�.b�������I�D%��#!}���qv\�%Yr;�񚢬o�<�|z!��mS�<A�����:�~���E����>`�;��60R}��f��g��׽WP4C*��A i��z���:��_��,��ar�Q�-��3�<�gl��BV`�I�`2X�iC�e���+�Dd���Nm�� ��n~��U��āC��	�S��6��40\���FW����J.NN{�����tFr,�4��@g�Xk���n��bnR�c�����w~r��C'�y�<�4�wC-�٭u�,*�^ �0�N���}\������~s��|uB��.6A��p�z�mw5��� ������Gl�R�ϸh���G��v��34uql��՚�Ǔ**�m`�i�B� ���¿g�I�o�x�������%!Z�xm%�t�=�8(��|L��e$�Ч��Wt�Q�����S'$�ց��$J��z�^6*+���VQ����R��a�h�CCZi�����p�����i��O�Pt�D�����(������6D����+������jY�4�6��S�A��X`���ֳGWہ�.�Y�;�j�+|q���£�M�x`IS��z<줔=5��ҡ�aj��^�y k���w
���[쯴��Z�Kk�G��=�%{�O�v-c�@�?�}��i���E\tc#�x�^��
"QU2��&'æ����U_֘y�T��Js��;����o��]	��p����'q\j��Y�z�	��Al�Լ��Xh
۾v "E	����lNuk|���:1lc`Щ��H�ח5�@Ĕڜ�0��
u[��bu|�O�~����Py�	b_�����j��f��>%߬��/
����Q�8y���_�f-�R��lA�R�}�R,#��Q���ݙ�5���קCF�K8&&�Qio٣��Ey̶.��\�������+��P<'	��%t$-�	����Ut31Ԧ���I*��&3���:�^w���R�uk{  ���?ת ce��U�r�BK�X�+�E ~��7ݫ�A�'���y�k!�#��CwI#��;@a���zK�`P�8�0?Co����L��l��m@P�&P�ghVI���_�v�}�������E(�����6:����Ww���}Ï�6��Vަ��qڍ��i�˹A�� jbN��l��jW����>��M5��L�O�